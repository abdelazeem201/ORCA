#######################################################################
####                                                               ####
####  The data contained in the file is created for educational    #### 
####  and training purposes only and are not recommended           ####
####  for fabrication                                              ####
####                                                               ####
#######################################################################
####                                                               ####
####  Copyright (C) 2013 Synopsys, Inc.                            ####
####                                                               ####
#######################################################################
####                                                               ####
####  The 32/28nm Generic Library ("Library") is unsupported       ####    
####  Confidential Information of Synopsys, Inc. ("Synopsys")      ####    
####  provided to you as Documentation under the terms of the      ####    
####  End User Software License Agreement between you or your      ####    
####  employer and Synopsys ("License Agreement") and you agree    ####    
####  not to distribute or disclose the Library without the        ####    
####  prior written consent of Synopsys. The Library IS NOT an     ####    
####  item of Licensed Software or Licensed Product under the      ####    
####  License Agreement.  Synopsys and/or its licensors own        ####    
####  and shall retain all right, title and interest in and        ####    
####  to the Library and all modifications thereto, including      ####    
####  all intellectual property rights embodied therein. All       ####    
####  rights in and to any Library modifications you make are      ####    
####  hereby assigned to Synopsys. If you do not agree with        ####    
####  this notice, including the disclaimer below, then you        ####    
####  are not authorized to use the Library.                       ####    
####                                                               ####  
####                                                               ####      
####  THIS LIBRARY IS BEING DISTRIBUTED BY SYNOPSYS SOLELY ON AN   ####
####  "AS IS" BASIS, WITH NO INTELLECUTAL PROPERTY                 ####
####  INDEMNIFICATION AND NO SUPPORT. ANY EXPRESS OR IMPLIED       ####
####  WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED       ####
####  WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR   ####
####  PURPOSE ARE HEREBY DISCLAIMED. IN NO EVENT SHALL SYNOPSYS    ####
####  BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     ####
####  EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT      ####
####  LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;     ####
####  LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)     ####
####  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN    ####
####  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE    ####
####  OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS      ####
####  DOCUMENTATION, EVEN IF ADVISED OF THE POSSIBILITY OF         ####
####  SUCH DAMAGE.                                                 #### 
####                                                               ####  
#######################################################################

# 
# LEF OUT 
# User Name : edbab 
# Date : Mon Dec 24 17:38:58 2012
# 
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "_<>" ;
DIVIDERCHAR "/" ;

MACRO SRAMLP1RW128x48
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 88.16 BY 238.887 ;
  SYMMETRY X Y R90 ;

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9600 17.2900 88.1600 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9600 17.2900 88.1600 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9600 17.2900 88.1600 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9600 17.2900 88.1600 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9600 17.2900 88.1600 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9600 16.8300 88.1600 17.0300 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9600 16.8300 88.1600 17.0300 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9600 16.8300 88.1600 17.0300 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9600 16.8300 88.1600 17.0300 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9600 16.8300 88.1600 17.0300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9600 9.8210 88.1600 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9600 9.8210 88.1600 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9600 9.8210 88.1600 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9600 9.8210 88.1600 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9600 9.8210 88.1600 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.4430 0.0000 21.6430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.4430 0.0000 21.6430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.4430 0.0000 21.6430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.4430 0.0000 21.6430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.4430 0.0000 21.6430 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[47]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1230 0.0000 35.3230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1230 0.0000 35.3230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1230 0.0000 35.3230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1230 0.0000 35.3230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1230 0.0000 35.3230 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[1]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3820 0.0000 45.5820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3820 0.0000 45.5820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3820 0.0000 45.5820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3820 0.0000 45.5820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3820 0.0000 45.5820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9740 0.0010 3.1740 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9740 0.0010 3.1740 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6590 0.0000 3.8590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6590 0.0000 3.8590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6590 0.0000 3.8590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6590 0.0000 3.8590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6590 0.0000 3.8590 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[21]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.0750 0.0000 20.2750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.0750 0.0000 20.2750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.0750 0.0000 20.2750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.0750 0.0000 20.2750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.0750 0.0000 20.2750 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[24]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9610 185.5460 88.1600 185.7460 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9610 185.5460 88.1600 185.7460 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9610 185.5460 88.1600 185.7460 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9610 185.5460 88.1600 185.7460 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9610 185.5460 88.1600 185.7460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9760 192.7680 88.1600 192.9680 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9760 192.7680 88.1600 192.9680 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9760 192.7680 88.1600 192.9680 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9760 192.7680 88.1600 192.9680 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9760 192.7680 88.1600 192.9680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9600 201.5900 88.1600 201.7900 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9600 201.5900 88.1600 201.7900 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9600 201.5900 88.1600 201.7900 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9600 201.5900 88.1600 201.7900 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9600 201.5900 88.1600 201.7900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9630 194.3660 88.1600 194.5660 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9630 194.3660 88.1600 194.5660 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9630 194.3660 88.1600 194.5660 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9630 194.3660 88.1600 194.5660 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9630 194.3660 88.1600 194.5660 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 84.9120 238.5870 85.2130 238.8870 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.8120 238.5870 86.1130 238.8870 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.0120 238.5870 84.3130 238.8870 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 35.8640 238.5860 36.1630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.0640 238.5860 34.3640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.9640 238.5860 35.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.3640 238.5860 40.6640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.0630 238.5860 43.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.5630 238.5860 38.8630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.2630 238.5860 41.5620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.4630 238.5860 39.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.6640 238.5860 46.9650 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.1640 238.5860 51.4650 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.7630 238.5860 46.0620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.9630 238.5860 44.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.5630 238.5860 47.8630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.2630 238.5860 50.5620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.3640 238.5860 49.6640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.4630 238.5860 48.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.8640 238.5860 45.1640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.4620 238.5860 57.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.6630 238.5860 1.9640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.0620 238.5860 61.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.2630 238.5860 5.5640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.8640 238.5860 54.1640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.0630 238.5860 52.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.6630 238.5860 55.9630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.7630 238.5860 55.0630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.9630 238.5860 53.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.2630 238.5860 59.5630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.4640 238.5860 3.7640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.3620 238.5860 58.6620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.5630 238.5860 2.8630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.5630 238.5860 56.8620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.7640 238.5860 1.0630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.1620 238.5860 60.4620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.3630 238.5860 4.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.5620 238.5860 65.8630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.7630 238.5860 10.0640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.4620 238.5860 66.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.6630 238.5860 10.9640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.9620 238.5860 62.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.1630 238.5860 6.4640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.6630 238.5860 64.9620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.8640 238.5860 9.1630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.3630 238.5860 67.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.5640 238.5860 11.8640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.1620 238.5860 69.4620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.3630 238.5860 13.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.7630 238.5860 64.0620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.9640 238.5860 8.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.8630 238.5860 63.1630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.0640 238.5860 7.3640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.2630 238.5860 68.5620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.4640 238.5860 12.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.6620 238.5860 73.9630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.8630 238.5860 18.1640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.4620 238.5860 75.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.6630 238.5860 19.9640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.5620 238.5860 74.8630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.7630 238.5860 19.0640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.3630 238.5860 76.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.5640 238.5860 20.8640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.7620 238.5860 73.0620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.9630 238.5860 17.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.8630 238.5860 72.1620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.0640 238.5860 16.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.0630 238.5860 70.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.2640 238.5860 14.5640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.9620 238.5860 71.2620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.1630 238.5860 15.4630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.7620 238.5860 82.0630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.9630 238.5860 26.2640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.0620 238.5860 79.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.2630 238.5860 23.5640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.4620 238.5860 84.7620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.6630 238.5860 28.9630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.6620 238.5860 82.9620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.8630 238.5860 27.1630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.5630 238.5860 83.8630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.7640 238.5860 28.0640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.2630 238.5860 86.5630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.3630 238.5860 85.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.5640 238.5860 29.8640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.9630 238.5860 80.2630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.1640 238.5860 24.4640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.1620 238.5860 78.4620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.3630 238.5860 22.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.8630 238.5860 81.1620 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.0640 238.5860 25.3630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.2630 238.5860 77.5630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.4640 238.5860 21.7640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.1640 238.5860 42.4650 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.1630 238.5860 33.4640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.6630 238.5860 37.9640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.7630 238.5860 37.0640 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.4640 238.5860 30.7630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.3640 238.5860 31.6630 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.2630 238.5860 32.5640 238.8860 ;
    END
  END VSS

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8110 0.0000 23.0110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8110 0.0000 23.0110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8110 0.0000 23.0110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8110 0.0000 23.0110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8110 0.0000 23.0110 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[45]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.5470 0.0000 25.7470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.5470 0.0000 25.7470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.5470 0.0000 25.7470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.5470 0.0000 25.7470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.5470 0.0000 25.7470 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[28]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9150 0.0000 27.1150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9150 0.0000 27.1150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9150 0.0000 27.1150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9150 0.0000 27.1150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9150 0.0000 27.1150 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[35]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.2830 0.0000 28.4830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.2830 0.0000 28.4830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.2830 0.0000 28.4830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.2830 0.0000 28.4830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.2830 0.0000 28.4830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[26]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.6510 0.0000 29.8510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.6510 0.0000 29.8510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.6510 0.0000 29.8510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.6510 0.0000 29.8510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.6510 0.0000 29.8510 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[19]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.3870 0.0000 32.5870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.3870 0.0000 32.5870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.3870 0.0000 32.5870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.3870 0.0000 32.5870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.3870 0.0000 32.5870 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[27]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.7550 0.0000 33.9550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.7550 0.0000 33.9550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.7550 0.0000 33.9550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.7550 0.0000 33.9550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.7550 0.0000 33.9550 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[25]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.8590 0.0000 38.0590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.8590 0.0000 38.0590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.8590 0.0000 38.0590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.8590 0.0000 38.0590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.8590 0.0000 38.0590 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[3]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.7470 0.0000 59.9470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.7470 0.0000 59.9470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.7470 0.0000 59.9470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.7470 0.0000 59.9470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.7470 0.0000 59.9470 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[16]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1150 0.0000 61.3150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1150 0.0000 61.3150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1150 0.0000 61.3150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1150 0.0000 61.3150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1150 0.0000 61.3150 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[17]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.4830 0.0000 62.6830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.4830 0.0000 62.6830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.4830 0.0000 62.6830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.4830 0.0000 62.6830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.4830 0.0000 62.6830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[18]

  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.8510 0.0000 64.0510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.8510 0.0000 64.0510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.8510 0.0000 64.0510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.8510 0.0000 64.0510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.8510 0.0000 64.0510 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[46]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2190 0.0000 65.4190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2190 0.0000 65.4190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2190 0.0000 65.4190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2190 0.0000 65.4190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2190 0.0000 65.4190 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[38]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.5870 0.0000 66.7870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.5870 0.0000 66.7870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.5870 0.0000 66.7870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.5870 0.0000 66.7870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.5870 0.0000 66.7870 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[36]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0270 0.0000 5.2270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0270 0.0000 5.2270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0270 0.0000 5.2270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0270 0.0000 5.2270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0270 0.0000 5.2270 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[9]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9630 176.7270 88.1600 176.9270 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9630 176.7270 88.1600 176.9270 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9630 176.7270 88.1600 176.9270 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9630 176.7270 88.1600 176.9270 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9630 176.7270 88.1600 176.9270 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9600 175.1280 88.1600 175.3280 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9600 175.1280 88.1600 175.3280 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9600 175.1280 88.1600 175.3280 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9600 175.1280 88.1600 175.3280 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9600 175.1280 88.1600 175.3280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9630 183.9500 88.1600 184.1500 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9630 183.9500 88.1600 184.1500 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9630 183.9500 88.1600 184.1500 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9630 183.9500 88.1600 184.1500 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9630 183.9500 88.1600 184.1500 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3310 0.0000 43.5310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3310 0.0000 43.5310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3310 0.0000 43.5310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3310 0.0000 43.5310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3310 0.0000 43.5310 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[41]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7500 0.0000 46.9500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7500 0.0000 46.9500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7500 0.0000 46.9500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7500 0.0000 46.9500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7500 0.0000 46.9500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[42]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1180 0.0000 48.3180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1180 0.0000 48.3180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1180 0.0000 48.3180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1180 0.0000 48.3180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1180 0.0000 48.3180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.4860 0.0000 49.6860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.4860 0.0000 49.6860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.4860 0.0000 49.6860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.4860 0.0000 49.6860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.4860 0.0000 49.6860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8540 0.0000 51.0540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8540 0.0000 51.0540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8540 0.0000 51.0540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8540 0.0000 51.0540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8540 0.0000 51.0540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2220 0.0000 52.4220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2220 0.0000 52.4220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2220 0.0000 52.4220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2220 0.0000 52.4220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2220 0.0000 52.4220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.5900 0.0000 53.7900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.5900 0.0000 53.7900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.5900 0.0000 53.7900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.5900 0.0000 53.7900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.5900 0.0000 53.7900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9580 0.0000 55.1580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9580 0.0000 55.1580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9580 0.0000 55.1580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9580 0.0000 55.1580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9580 0.0000 55.1580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3260 0.0000 56.5260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3260 0.0000 56.5260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3260 0.0000 56.5260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3260 0.0000 56.5260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3260 0.0000 56.5260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.6940 0.0000 57.8940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.6940 0.0000 57.8940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.6940 0.0000 57.8940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.6940 0.0000 57.8940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.6940 0.0000 57.8940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0620 0.0000 59.2620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0620 0.0000 59.2620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0620 0.0000 59.2620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0620 0.0000 59.2620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0620 0.0000 59.2620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4300 0.0000 60.6300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4300 0.0000 60.6300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4300 0.0000 60.6300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4300 0.0000 60.6300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4300 0.0000 60.6300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.7980 0.0000 61.9980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.7980 0.0000 61.9980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.7980 0.0000 61.9980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.7980 0.0000 61.9980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.7980 0.0000 61.9980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1660 0.0000 63.3660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1660 0.0000 63.3660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1660 0.0000 63.3660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1660 0.0000 63.3660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1660 0.0000 63.3660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[46]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5340 0.0000 64.7340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5340 0.0000 64.7340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5340 0.0000 64.7340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5340 0.0000 64.7340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5340 0.0000 64.7340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.9020 0.0000 66.1020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.9020 0.0000 66.1020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.9020 0.0000 66.1020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.9020 0.0000 66.1020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.9020 0.0000 66.1020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.2600 0.0000 67.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.2600 0.0000 67.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.2600 0.0000 67.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.2600 0.0000 67.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.2600 0.0000 67.4600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2910 0.0000 2.4910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2910 0.0000 2.4910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2910 0.0000 2.4910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2910 0.0000 2.4910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2910 0.0000 2.4910 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[44]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.4990 0.0000 10.6990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.4990 0.0000 10.6990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.4990 0.0000 10.6990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.4990 0.0000 10.6990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.4990 0.0000 10.6990 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[39]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7630 0.0000 7.9630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7630 0.0000 7.9630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7630 0.0000 7.9630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7630 0.0000 7.9630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7630 0.0000 7.9630 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[11]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8030 0.0000 49.0030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8030 0.0000 49.0030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8030 0.0000 49.0030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8030 0.0000 49.0030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8030 0.0000 49.0030 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[7]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1740 0.0000 37.3740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1740 0.0000 37.3740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1740 0.0000 37.3740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1740 0.0000 37.3740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1740 0.0000 37.3740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4380 0.0000 34.6380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4380 0.0000 34.6380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4380 0.0000 34.6380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4380 0.0000 34.6380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4380 0.0000 34.6380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.9630 0.0000 42.1630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.9630 0.0000 42.1630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.9630 0.0000 42.1630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.9630 0.0000 42.1630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.9630 0.0000 42.1630 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[5]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0190 0.0000 31.2190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0190 0.0000 31.2190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0190 0.0000 31.2190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0190 0.0000 31.2190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0190 0.0000 31.2190 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[13]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7020 0.0000 31.9020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7020 0.0000 31.9020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7020 0.0000 31.9020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7020 0.0000 31.9020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7020 0.0000 31.9020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.1790 0.0000 24.3790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.1790 0.0000 24.3790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.1790 0.0000 24.3790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.1790 0.0000 24.3790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.1790 0.0000 24.3790 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[0]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8620 0.0000 25.0620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8620 0.0000 25.0620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8620 0.0000 25.0620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8620 0.0000 25.0620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8620 0.0000 25.0620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5950 0.0000 40.7950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5950 0.0000 40.7950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5950 0.0000 40.7950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5950 0.0000 40.7950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5950 0.0000 40.7950 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[40]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.0670 0.0000 46.2670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.0670 0.0000 46.2670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.0670 0.0000 46.2670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.0670 0.0000 46.2670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.0670 0.0000 46.2670 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[30]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0140 0.0000 44.2140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0140 0.0000 44.2140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0140 0.0000 44.2140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0140 0.0000 44.2140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0140 0.0000 44.2140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1310 0.0000 9.3310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1310 0.0000 9.3310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1310 0.0000 9.3310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1310 0.0000 9.3310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1310 0.0000 9.3310 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[10]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[39]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8060 0.0000 36.0060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8060 0.0000 36.0060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8060 0.0000 36.0060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8060 0.0000 36.0060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8060 0.0000 36.0060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2780 0.0000 41.4780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2780 0.0000 41.4780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2780 0.0000 41.4780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2780 0.0000 41.4780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2780 0.0000 41.4780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 19.3900 0.0000 19.5900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.3900 0.0000 19.5900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.3900 0.0000 19.5900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.3900 0.0000 19.5900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 19.3900 0.0000 19.5900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.1710 0.0000 50.3710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.1710 0.0000 50.3710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.1710 0.0000 50.3710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.1710 0.0000 50.3710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.1710 0.0000 50.3710 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[31]

  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.7580 0.0000 20.9580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.7580 0.0000 20.9580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.7580 0.0000 20.9580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.7580 0.0000 20.9580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.7580 0.0000 20.9580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[47]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9070 0.0000 53.1070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9070 0.0000 53.1070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9070 0.0000 53.1070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9070 0.0000 53.1070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9070 0.0000 53.1070 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[20]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5390 0.0000 51.7390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5390 0.0000 51.7390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5390 0.0000 51.7390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5390 0.0000 51.7390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5390 0.0000 51.7390 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[43]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.1260 0.0000 22.3260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.1260 0.0000 22.3260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.1260 0.0000 22.3260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.1260 0.0000 22.3260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.1260 0.0000 22.3260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4940 0.0000 23.6940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4940 0.0000 23.6940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4940 0.0000 23.6940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4940 0.0000 23.6940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4940 0.0000 23.6940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.2750 0.0000 54.4750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.2750 0.0000 54.4750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.2750 0.0000 54.4750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.2750 0.0000 54.4750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.2750 0.0000 54.4750 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[8]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0700 0.0000 33.2700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0700 0.0000 33.2700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0700 0.0000 33.2700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0700 0.0000 33.2700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0700 0.0000 33.2700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.6990 0.0000 44.8990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.6990 0.0000 44.8990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.6990 0.0000 44.8990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.6990 0.0000 44.8990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.6990 0.0000 44.8990 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[6]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2300 0.0000 26.4300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2300 0.0000 26.4300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2300 0.0000 26.4300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2300 0.0000 26.4300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2300 0.0000 26.4300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0110 0.0000 57.2110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0110 0.0000 57.2110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0110 0.0000 57.2110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0110 0.0000 57.2110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0110 0.0000 57.2110 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[14]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9660 0.0000 29.1660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9660 0.0000 29.1660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9660 0.0000 29.1660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9660 0.0000 29.1660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9660 0.0000 29.1660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.5980 0.0000 27.7980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.5980 0.0000 27.7980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.5980 0.0000 27.7980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.5980 0.0000 27.7980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.5980 0.0000 27.7980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4910 0.0000 36.6910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4910 0.0000 36.6910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4910 0.0000 36.6910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4910 0.0000 36.6910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4910 0.0000 36.6910 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[2]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2270 0.0000 39.4270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2270 0.0000 39.4270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2270 0.0000 39.4270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2270 0.0000 39.4270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2270 0.0000 39.4270 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[4]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3340 0.0000 30.5340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3340 0.0000 30.5340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3340 0.0000 30.5340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3340 0.0000 30.5340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3340 0.0000 30.5340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3950 0.0000 6.5950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3950 0.0000 6.5950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3950 0.0000 6.5950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3950 0.0000 6.5950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3950 0.0000 6.5950 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[12]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.7070 0.0000 18.9070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.7070 0.0000 18.9070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.7070 0.0000 18.9070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.7070 0.0000 18.9070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.7070 0.0000 18.9070 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[23]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6460 0.0000 42.8460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6460 0.0000 42.8460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6460 0.0000 42.8460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6460 0.0000 42.8460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6460 0.0000 42.8460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[41]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 17.3390 0.0000 17.5390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.3390 0.0000 17.5390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.3390 0.0000 17.5390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 17.3390 0.0000 17.5390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 17.3390 0.0000 17.5390 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[29]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9100 0.0000 40.1100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9100 0.0000 40.1100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9100 0.0000 40.1100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9100 0.0000 40.1100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9100 0.0000 40.1100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[40]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5420 0.0000 38.7420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5420 0.0000 38.7420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5420 0.0000 38.7420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5420 0.0000 38.7420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5420 0.0000 38.7420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.9710 0.0000 16.1710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.9710 0.0000 16.1710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.9710 0.0000 16.1710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.9710 0.0000 16.1710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.9710 0.0000 16.1710 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[33]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[37]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.2350 0.0000 13.4350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.2350 0.0000 13.4350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.2350 0.0000 13.4350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.2350 0.0000 13.4350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.2350 0.0000 13.4350 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[34]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8670 0.0000 12.0670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8670 0.0000 12.0670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8670 0.0000 12.0670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8670 0.0000 12.0670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8670 0.0000 12.0670 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[37]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.6030 0.0000 14.8030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.6030 0.0000 14.8030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.6030 0.0000 14.8030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.6030 0.0000 14.8030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.6030 0.0000 14.8030 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[22]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.2860 0.0000 15.4860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.2860 0.0000 15.4860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.2860 0.0000 15.4860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.2860 0.0000 15.4860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.2860 0.0000 15.4860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.9180 0.0000 14.1180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.9180 0.0000 14.1180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.9180 0.0000 14.1180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.9180 0.0000 14.1180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.9180 0.0000 14.1180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.3790 0.0000 58.5790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.3790 0.0000 58.5790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.3790 0.0000 58.5790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.3790 0.0000 58.5790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.3790 0.0000 58.5790 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[15]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.6540 0.0000 16.8540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.6540 0.0000 16.8540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.6540 0.0000 16.8540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.6540 0.0000 16.8540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.6540 0.0000 16.8540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4350 0.0000 47.6350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4350 0.0000 47.6350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4350 0.0000 47.6350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4350 0.0000 47.6350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4350 0.0000 47.6350 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[42]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.0220 0.0000 18.2220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.0220 0.0000 18.2220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.0220 0.0000 18.2220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.0220 0.0000 18.2220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.0220 0.0000 18.2220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.6430 0.0000 55.8430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.6430 0.0000 55.8430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.6430 0.0000 55.8430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.6430 0.0000 55.8430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.6430 0.0000 55.8430 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[32]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.0130 238.5860 75.3130 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.9120 238.5860 76.2130 238.8860 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.8130 238.5860 77.1130 238.8860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9660 221.3070 88.1600 221.5070 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9660 221.3070 88.1600 221.5070 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9660 221.3070 88.1600 221.5070 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9660 221.3070 88.1600 221.5070 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9660 221.3070 88.1600 221.5070 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9660 218.0550 88.1600 218.2550 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9660 218.0550 88.1600 218.2550 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9660 218.0550 88.1600 218.2550 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9660 218.0550 88.1600 218.2550 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9660 218.0550 88.1600 218.2550 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9660 217.7120 88.1600 217.9120 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9660 217.7120 88.1600 217.9120 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9660 217.7120 88.1600 217.9120 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9660 217.7120 88.1600 217.9120 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9660 217.7120 88.1600 217.9120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD
  OBS
    LAYER M2 ;
      RECT 0.0000 174.4280 87.2600 176.0280 ;
      RECT 0.0000 18.1900 88.1600 174.4280 ;
      RECT 0.0000 16.1300 87.2600 18.1900 ;
      RECT 0.0000 10.7210 88.1600 16.1300 ;
      RECT 0.0000 9.1210 87.2600 10.7210 ;
      RECT 0.0000 0.9000 88.1600 9.1210 ;
      RECT 68.1600 0.0000 88.1600 9.1210 ;
      RECT 68.1600 0.0000 88.1600 0.9000 ;
      RECT 0.0000 222.2070 88.1600 238.8870 ;
      RECT 0.0000 202.4900 87.2660 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 217.0120 87.2660 222.2070 ;
      RECT 0.0000 202.4900 88.1600 217.0120 ;
      RECT 0.0000 200.8900 87.2600 202.4900 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 86.6590 218.9550 88.1600 220.6070 ;
      RECT 0.0000 195.2660 88.1600 200.8900 ;
      RECT 0.0000 186.4460 87.2630 200.8900 ;
      RECT 0.0000 176.0280 87.2610 200.8900 ;
      RECT 0.0000 193.6660 87.2630 195.2660 ;
      RECT 0.0000 192.0680 87.2760 193.6660 ;
      RECT 0.0000 186.4460 87.2760 193.6660 ;
      RECT 0.0000 186.4460 88.1600 192.0680 ;
      RECT 0.0000 184.8460 87.2610 186.4460 ;
      RECT 0.0000 183.2500 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 177.6270 88.1600 183.2500 ;
      RECT 0.0000 176.0280 87.2630 177.6270 ;
    LAYER M1 ;
      RECT 87.3630 175.9280 88.1600 176.1270 ;
      RECT 87.3760 193.5680 88.1600 193.7660 ;
      RECT 87.3630 184.7500 88.1600 184.9460 ;
      RECT 0.0000 0.0000 1.0060 0.8000 ;
      RECT 86.6590 218.8550 88.1600 220.7070 ;
      RECT 0.0000 195.1660 88.1600 200.9900 ;
      RECT 0.0000 186.3460 87.3630 200.9900 ;
      RECT 0.0000 175.9280 87.3610 200.9900 ;
      RECT 0.0000 193.7660 87.3630 195.1660 ;
      RECT 0.0000 192.1680 87.3760 193.7660 ;
      RECT 0.0000 186.3460 87.3760 193.7660 ;
      RECT 0.0000 186.3460 88.1600 192.1680 ;
      RECT 0.0000 184.9460 87.3610 186.3460 ;
      RECT 0.0000 183.3500 87.3630 184.9460 ;
      RECT 0.0000 175.9280 87.3630 184.9460 ;
      RECT 0.0000 175.9280 87.3630 184.9460 ;
      RECT 0.0000 177.5270 88.1600 183.3500 ;
      RECT 0.0000 175.9280 87.3630 177.5270 ;
      RECT 0.0000 174.5280 87.3600 175.9280 ;
      RECT 0.0000 18.0900 88.1600 174.5280 ;
      RECT 0.0000 16.2300 87.3600 18.0900 ;
      RECT 0.0000 10.6210 88.1600 16.2300 ;
      RECT 0.0000 9.2210 87.3600 10.6210 ;
      RECT 0.0000 0.8000 88.1600 9.2210 ;
      RECT 68.0600 0.0000 88.1600 9.2210 ;
      RECT 68.0600 0.0000 88.1600 0.8000 ;
      RECT 0.0000 222.1070 88.1600 238.8870 ;
      RECT 0.0000 202.3900 87.3660 238.8870 ;
      RECT 0.0000 0.8000 87.3600 238.8870 ;
      RECT 0.0000 0.8000 87.3600 238.8870 ;
      RECT 0.0000 0.8000 87.3600 238.8870 ;
      RECT 0.0000 0.8000 87.3600 238.8870 ;
      RECT 0.0000 217.1120 87.3660 222.1070 ;
      RECT 0.0000 202.3900 88.1600 217.1120 ;
      RECT 0.0000 200.9900 87.3600 202.3900 ;
    LAYER PO ;
      RECT 0.0000 0.0000 88.1600 238.8870 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 88.1600 238.8870 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 88.1600 238.8870 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 88.1600 238.8870 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 88.1600 238.8870 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 88.1600 238.8870 ;
    LAYER M5 ;
      RECT 0.0000 237.8860 0.0640 238.8870 ;
      RECT 0.0000 0.0000 0.9060 0.9010 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 87.2630 237.8860 88.1600 238.8870 ;
      RECT 0.0000 0.9000 2.2740 0.9010 ;
      RECT 0.0000 0.9000 2.2740 2.4010 ;
      RECT 86.6590 218.9550 88.1600 220.6070 ;
      RECT 68.1600 0.0000 88.1600 0.9000 ;
      RECT 0.0000 195.2660 88.1600 200.8900 ;
      RECT 0.0000 186.4460 87.2630 200.8900 ;
      RECT 0.0000 176.0280 87.2610 200.8900 ;
      RECT 0.0000 193.6660 87.2630 195.2660 ;
      RECT 0.0000 192.0680 87.2760 193.6660 ;
      RECT 0.0000 186.4460 87.2760 193.6660 ;
      RECT 0.0000 186.4460 88.1600 192.0680 ;
      RECT 0.0000 184.8460 87.2610 186.4460 ;
      RECT 0.0000 183.2500 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 177.6270 88.1600 183.2500 ;
      RECT 0.0000 176.0280 87.2630 177.6270 ;
      RECT 0.0000 174.4280 87.2600 176.0280 ;
      RECT 0.0000 18.1900 88.1600 174.4280 ;
      RECT 0.0000 16.1300 87.2600 18.1900 ;
      RECT 0.0000 10.7210 88.1600 16.1300 ;
      RECT 0.0000 9.1210 87.2600 10.7210 ;
      RECT 0.0000 0.9010 88.1600 9.1210 ;
      RECT 3.8740 0.9000 88.1600 9.1210 ;
      RECT 3.8740 0.9000 88.1600 0.9010 ;
      RECT 68.1600 0.0000 88.1600 9.1210 ;
      RECT 0.0000 222.2070 88.1600 237.8860 ;
      RECT 0.0000 202.4900 87.2660 237.8860 ;
      RECT 0.0000 0.9010 87.2600 237.8860 ;
      RECT 0.0000 0.9010 87.2600 237.8860 ;
      RECT 0.0000 0.9010 87.2600 237.8860 ;
      RECT 0.0000 0.9010 87.2600 237.8860 ;
      RECT 0.0000 217.0120 87.2660 222.2070 ;
      RECT 0.0000 202.4900 88.1600 217.0120 ;
      RECT 0.0000 200.8900 87.2600 202.4900 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9060 0.9010 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 0.0000 0.9000 2.2740 2.4010 ;
      RECT 86.6590 218.9550 88.1600 220.6070 ;
      RECT 68.1600 0.0000 88.1600 0.9000 ;
      RECT 0.0000 195.2660 88.1600 200.8900 ;
      RECT 0.0000 186.4460 87.2630 200.8900 ;
      RECT 0.0000 176.0280 87.2610 200.8900 ;
      RECT 0.0000 193.6660 87.2630 195.2660 ;
      RECT 0.0000 192.0680 87.2760 193.6660 ;
      RECT 0.0000 186.4460 87.2760 193.6660 ;
      RECT 0.0000 186.4460 88.1600 192.0680 ;
      RECT 0.0000 184.8460 87.2610 186.4460 ;
      RECT 0.0000 183.2500 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 177.6270 88.1600 183.2500 ;
      RECT 0.0000 176.0280 87.2630 177.6270 ;
      RECT 0.0000 174.4280 87.2600 176.0280 ;
      RECT 0.0000 18.1900 88.1600 174.4280 ;
      RECT 0.0000 16.1300 87.2600 18.1900 ;
      RECT 0.0000 10.7210 88.1600 16.1300 ;
      RECT 0.0000 9.1210 87.2600 10.7210 ;
      RECT 0.0000 0.9010 88.1600 9.1210 ;
      RECT 3.8740 0.9000 88.1600 9.1210 ;
      RECT 3.8740 0.9000 88.1600 0.9010 ;
      RECT 68.1600 0.0000 88.1600 9.1210 ;
      RECT 0.0000 222.2070 88.1600 238.8870 ;
      RECT 0.0000 202.4900 87.2660 238.8870 ;
      RECT 0.0000 0.9010 87.2600 238.8870 ;
      RECT 0.0000 0.9010 87.2600 238.8870 ;
      RECT 0.0000 0.9010 87.2600 238.8870 ;
      RECT 0.0000 0.9010 87.2600 238.8870 ;
      RECT 0.0000 217.0120 87.2660 222.2070 ;
      RECT 0.0000 202.4900 88.1600 217.0120 ;
      RECT 0.0000 200.8900 87.2600 202.4900 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 86.6590 218.9550 88.1600 220.6070 ;
      RECT 0.0000 195.2660 88.1600 200.8900 ;
      RECT 0.0000 186.4460 87.2630 200.8900 ;
      RECT 0.0000 176.0280 87.2610 200.8900 ;
      RECT 0.0000 193.6660 87.2630 195.2660 ;
      RECT 0.0000 192.0680 87.2760 193.6660 ;
      RECT 0.0000 186.4460 87.2760 193.6660 ;
      RECT 0.0000 186.4460 88.1600 192.0680 ;
      RECT 0.0000 184.8460 87.2610 186.4460 ;
      RECT 0.0000 183.2500 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 176.0280 87.2630 184.8460 ;
      RECT 0.0000 177.6270 88.1600 183.2500 ;
      RECT 0.0000 176.0280 87.2630 177.6270 ;
      RECT 0.0000 174.4280 87.2600 176.0280 ;
      RECT 0.0000 18.1900 88.1600 174.4280 ;
      RECT 0.0000 16.1300 87.2600 18.1900 ;
      RECT 0.0000 10.7210 88.1600 16.1300 ;
      RECT 0.0000 9.1210 87.2600 10.7210 ;
      RECT 0.0000 0.9000 88.1600 9.1210 ;
      RECT 68.1600 0.0000 88.1600 9.1210 ;
      RECT 68.1600 0.0000 88.1600 0.9000 ;
      RECT 0.0000 222.2070 88.1600 238.8870 ;
      RECT 0.0000 202.4900 87.2660 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 0.9000 87.2600 238.8870 ;
      RECT 0.0000 217.0120 87.2660 222.2070 ;
      RECT 0.0000 202.4900 88.1600 217.0120 ;
      RECT 0.0000 200.8900 87.2600 202.4900 ;
  END
END SRAMLP1RW128x48

MACRO SRAMLP1RW256x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 38.137 BY 247.882 ;
  SYMMETRY X Y R90 ;

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9370 16.8970 38.1370 17.0970 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9370 16.8970 38.1370 17.0970 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9370 16.8970 38.1370 17.0970 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9370 16.8970 38.1370 17.0970 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9370 16.8970 38.1370 17.0970 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9370 180.8310 38.1370 181.0310 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9370 180.8310 38.1370 181.0310 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9370 180.8310 38.1370 181.0310 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9370 180.8310 38.1370 181.0310 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9370 180.8310 38.1370 181.0310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9400 182.4300 38.1370 182.6300 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9400 182.4300 38.1370 182.6300 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9400 182.4300 38.1370 182.6300 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9400 182.4300 38.1370 182.6300 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9400 182.4300 38.1370 182.6300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.6940 0.0000 4.8940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.6940 0.0000 4.8940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.6940 0.0000 4.8940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.6940 0.0000 4.8940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.6940 0.0000 4.8940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.9890 0.0000 4.1890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.9890 0.0000 4.1890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.9890 0.0000 4.1890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.9890 0.0000 4.1890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.9890 0.0000 4.1890 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[2]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.4640 0.0000 9.6640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.4640 0.0000 9.6640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.4640 0.0000 9.6640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.4640 0.0000 9.6640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.4640 0.0000 9.6640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[3]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.8340 0.0000 11.0340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.8340 0.0000 11.0340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.8340 0.0000 11.0340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.8340 0.0000 11.0340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.8340 0.0000 11.0340 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[4]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.1660 0.0000 10.3660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.1660 0.0000 10.3660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.1660 0.0000 10.3660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.1660 0.0000 10.3660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.1660 0.0000 10.3660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.3590 0.0000 5.5590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.3590 0.0000 5.5590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.3590 0.0000 5.5590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.3590 0.0000 5.5590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.3590 0.0000 5.5590 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[5]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.3260 0.0000 3.5260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.3260 0.0000 3.5260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.3260 0.0000 3.5260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.3260 0.0000 3.5260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.3260 0.0000 3.5260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9370 17.3630 38.1370 17.5630 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9370 17.3630 38.1370 17.5630 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9370 17.3630 38.1370 17.5630 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9370 17.3630 38.1370 17.5630 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9370 17.3630 38.1370 17.5630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9400 189.6530 38.1370 189.8530 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9400 189.6530 38.1370 189.8530 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9400 189.6530 38.1370 189.8530 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9400 189.6530 38.1370 189.8530 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9400 189.6530 38.1370 189.8530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9370 9.8900 38.1370 10.0900 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9370 9.8900 38.1370 10.0900 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9370 9.8900 38.1370 10.0900 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9370 9.8900 38.1370 10.0900 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9370 9.8900 38.1370 10.0900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9380 191.2490 38.1370 191.4490 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9380 191.2490 38.1370 191.4490 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9380 191.2490 38.1370 191.4490 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9380 191.2490 38.1370 191.4490 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9380 191.2490 38.1370 191.4490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.0820 0.0000 8.2820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.0820 0.0000 8.2820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.0820 0.0000 8.2820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.0820 0.0000 8.2820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.0820 0.0000 8.2820 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564528 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564528 LAYER M3 ;
  END O[7]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9400 200.0690 38.1370 200.2690 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9400 200.0690 38.1370 200.2690 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9400 200.0690 38.1370 200.2690 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9400 200.0690 38.1370 200.2690 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9400 200.0690 38.1370 200.2690 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9430 223.9160 38.1370 224.1160 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9430 223.9160 38.1370 224.1160 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9430 223.9160 38.1370 224.1160 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9430 223.9160 38.1370 224.1160 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9430 223.9160 38.1370 224.1160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9370 207.2930 38.1370 207.4930 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9370 207.2930 38.1370 207.4930 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9370 207.2930 38.1370 207.4930 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9370 207.2930 38.1370 207.4930 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9370 207.2930 38.1370 207.4930 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9430 227.4820 38.1370 227.6820 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9430 227.4820 38.1370 227.6820 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9430 227.4820 38.1370 227.6820 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9430 227.4820 38.1370 227.6820 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9430 227.4820 38.1370 227.6820 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9530 198.4710 38.1370 198.6710 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9530 198.4710 38.1370 198.6710 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9530 198.4710 38.1370 198.6710 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9530 198.4710 38.1370 198.6710 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9530 198.4710 38.1370 198.6710 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.5540 247.5760 26.8530 247.8780 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.4550 247.5760 27.7540 247.8780 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.3550 247.5760 28.6550 247.8780 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.9010 0.0000 13.1010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.9010 0.0000 13.1010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.9010 0.0000 13.1010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.9010 0.0000 13.1010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.9010 0.0000 13.1010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9370 29.3920 38.1370 29.5920 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9370 29.3920 38.1370 29.5920 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9370 29.3920 38.1370 29.5920 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9370 29.3920 38.1370 29.5920 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9370 29.3920 38.1370 29.5920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9430 224.2960 38.1370 224.4960 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9430 224.2960 38.1370 224.4960 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9430 224.2960 38.1370 224.4960 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9430 224.2960 38.1370 224.4960 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9430 224.2960 38.1370 224.4960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.4300 0.0000 7.6300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.4300 0.0000 7.6300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.4300 0.0000 7.6300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.4300 0.0000 7.6300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.4300 0.0000 7.6300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.7280 0.0000 6.9280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.7280 0.0000 6.9280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.7280 0.0000 6.9280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.7280 0.0000 6.9280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.7280 0.0000 6.9280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[6]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.0620 0.0000 6.2620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.0620 0.0000 6.2620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.0620 0.0000 6.2620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.0620 0.0000 6.2620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.0620 0.0000 6.2620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.2040 0.0000 12.4040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.2040 0.0000 12.4040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.2040 0.0000 12.4040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.2040 0.0000 12.4040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.2040 0.0000 12.4040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[0]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 34.6550 247.5760 34.9550 247.8780 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.5540 247.5760 35.8540 247.8780 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.4540 247.5760 36.7540 247.8780 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.5030 247.5800 4.8040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.4030 247.5800 14.7030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.8030 247.5800 11.1030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7040 247.5800 3.0030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.2040 247.5800 16.5040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1030 247.5800 17.4020 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.3030 247.5800 15.6030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0040 247.5800 18.3050 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.2040 247.5800 7.5040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7040 247.5800 12.0040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.5040 247.5800 13.8050 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6030 247.5800 12.9020 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.1030 247.5800 8.4020 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.9030 247.5800 10.2030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.0040 247.5800 9.3050 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.0030 247.5800 36.3030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.5030 247.5800 31.8030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.9040 247.5800 28.2040 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.3040 247.5800 24.6040 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.7040 247.5800 21.0040 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.9030 247.5800 19.2030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.9020 247.5800 37.2020 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.1020 247.5800 35.4020 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.2030 247.5800 34.5030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.3030 247.5800 33.6030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.4020 247.5800 32.7020 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.6020 247.5800 30.9020 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.7030 247.5800 30.0030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.8030 247.5800 29.1030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.0030 247.5800 27.3030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.1030 247.5800 26.4030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.2030 247.5800 25.5030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.4030 247.5800 23.7030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.5030 247.5800 22.8030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.6030 247.5800 21.9030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.8030 247.5800 20.1030 247.8820 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.8040 247.5800 2.1030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.9040 247.5800 1.2040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0040 247.5800 0.3040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.4030 247.5800 5.7030 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6030 247.5800 3.9040 247.8800 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.3030 247.5800 6.6030 247.8800 ;
    END
    ANTENNAPARTIALMETALAREA 74.03999 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 74.03999 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 74.0394 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 74.0394 LAYER M5 ;
  END VSS

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.6120 0.0000 2.8120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.6120 0.0000 2.8120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.6120 0.0000 2.8120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.6120 0.0000 2.8120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.6120 0.0000 2.8120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.564648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.564648 LAYER M3 ;
  END O[1]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.5340 0.0000 11.7340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.5340 0.0000 11.7340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.5340 0.0000 11.7340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.5340 0.0000 11.7340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.5340 0.0000 11.7340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.9580 0.0000 2.1580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.9580 0.0000 2.1580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.9580 0.0000 2.1580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.9580 0.0000 2.1580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.9580 0.0000 2.1580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.7980 0.0000 8.9980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.7980 0.0000 8.9980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.7980 0.0000 8.9980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.7980 0.0000 8.9980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.7980 0.0000 8.9980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]
  OBS
    LAYER M2 ;
      RECT 0.0000 188.9530 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 183.3300 38.1370 188.9530 ;
      RECT 0.0000 181.7310 37.2400 183.3300 ;
      RECT 0.0000 180.1310 37.2370 181.7310 ;
      RECT 0.0000 30.2920 38.1370 180.1310 ;
      RECT 0.0000 28.6920 37.2370 30.2920 ;
      RECT 0.0000 18.2630 38.1370 28.6920 ;
      RECT 0.0000 16.1970 37.2370 18.2630 ;
      RECT 0.0000 10.7900 38.1370 16.1970 ;
      RECT 0.0000 9.1900 37.2370 10.7900 ;
      RECT 0.0000 0.9000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 0.9000 ;
      RECT 0.0000 228.3820 38.1370 247.8820 ;
      RECT 0.0000 208.1930 37.2430 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 223.2160 37.2430 228.3820 ;
      RECT 0.0000 208.1930 38.1370 223.2160 ;
      RECT 0.0000 206.5930 37.2370 208.1930 ;
      RECT 0.0000 0.0000 1.2580 0.9000 ;
      RECT 36.6360 225.1960 38.1370 226.7820 ;
      RECT 0.0000 200.9690 38.1370 206.5930 ;
      RECT 0.0000 192.1490 37.2400 206.5930 ;
      RECT 0.0000 181.7310 37.2380 206.5930 ;
      RECT 0.0000 199.3690 37.2400 200.9690 ;
      RECT 0.0000 197.7710 37.2530 199.3690 ;
      RECT 0.0000 192.1490 37.2530 199.3690 ;
      RECT 0.0000 192.1490 38.1370 197.7710 ;
      RECT 0.0000 190.5490 37.2380 192.1490 ;
    LAYER M1 ;
      RECT 37.3400 190.4530 38.1370 190.6490 ;
      RECT 37.3530 199.2710 38.1370 199.4690 ;
      RECT 37.3400 181.6310 38.1370 181.8300 ;
      RECT 0.0000 0.0000 1.3580 0.8000 ;
      RECT 36.6360 225.0960 38.1370 226.8820 ;
      RECT 0.0000 200.8690 38.1370 206.6930 ;
      RECT 0.0000 192.0490 37.3400 206.6930 ;
      RECT 0.0000 181.6310 37.3380 206.6930 ;
      RECT 0.0000 199.4690 37.3400 200.8690 ;
      RECT 0.0000 197.8710 37.3530 199.4690 ;
      RECT 0.0000 192.0490 37.3530 199.4690 ;
      RECT 0.0000 192.0490 38.1370 197.8710 ;
      RECT 0.0000 190.6490 37.3380 192.0490 ;
      RECT 0.0000 189.0530 37.3400 190.6490 ;
      RECT 0.0000 181.6310 37.3400 190.6490 ;
      RECT 0.0000 181.6310 37.3400 190.6490 ;
      RECT 0.0000 183.2300 38.1370 189.0530 ;
      RECT 0.0000 181.6310 37.3400 183.2300 ;
      RECT 0.0000 180.2310 37.3370 181.6310 ;
      RECT 0.0000 30.1920 38.1370 180.2310 ;
      RECT 0.0000 28.7920 37.3370 30.1920 ;
      RECT 0.0000 18.1630 38.1370 28.7920 ;
      RECT 0.0000 16.2970 37.3370 18.1630 ;
      RECT 0.0000 10.6900 38.1370 16.2970 ;
      RECT 0.0000 9.2900 37.3370 10.6900 ;
      RECT 0.0000 0.8000 38.1370 9.2900 ;
      RECT 13.7010 0.0000 38.1370 9.2900 ;
      RECT 13.7010 0.0000 38.1370 0.8000 ;
      RECT 0.0000 228.2820 38.1370 247.8820 ;
      RECT 0.0000 208.0930 37.3430 247.8820 ;
      RECT 0.0000 0.8000 37.3370 247.8820 ;
      RECT 0.0000 0.8000 37.3370 247.8820 ;
      RECT 0.0000 0.8000 37.3370 247.8820 ;
      RECT 0.0000 0.8000 37.3370 247.8820 ;
      RECT 0.0000 0.8000 37.3370 247.8820 ;
      RECT 0.0000 223.3160 37.3430 228.2820 ;
      RECT 0.0000 208.0930 38.1370 223.3160 ;
      RECT 0.0000 206.6930 37.3370 208.0930 ;
    LAYER PO ;
      RECT 0.0000 0.0000 38.1370 247.8820 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 38.1370 247.8820 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 38.1370 247.8820 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 38.1370 247.8820 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 38.1370 247.8820 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 38.1370 247.8820 ;
    LAYER M5 ;
      RECT 37.9020 246.8800 38.1370 247.8820 ;
      RECT 0.0000 0.0000 1.2580 0.9000 ;
      RECT 37.4540 246.8760 38.1370 246.8800 ;
      RECT 36.6360 225.1960 38.1370 226.7820 ;
      RECT 37.4540 246.5790 38.1370 246.8800 ;
      RECT 0.0000 246.8760 25.8540 246.8800 ;
      RECT 0.0000 0.9000 25.8540 246.8800 ;
      RECT 0.0000 228.3820 38.1370 246.8760 ;
      RECT 0.0000 208.1930 37.2430 246.8760 ;
      RECT 0.0000 0.9000 37.2370 246.8760 ;
      RECT 0.0000 0.9000 37.2370 246.8760 ;
      RECT 0.0000 0.9000 37.2370 246.8760 ;
      RECT 0.0000 0.9000 37.2370 246.8760 ;
      RECT 0.0000 0.9000 37.2370 246.8760 ;
      RECT 0.0000 223.2160 37.2430 228.3820 ;
      RECT 0.0000 208.1930 38.1370 223.2160 ;
      RECT 0.0000 206.5930 37.2370 208.1930 ;
      RECT 0.0000 200.9690 38.1370 206.5930 ;
      RECT 0.0000 192.1490 37.2400 206.5930 ;
      RECT 0.0000 181.7310 37.2380 206.5930 ;
      RECT 0.0000 199.3690 37.2400 200.9690 ;
      RECT 0.0000 197.7710 37.2530 199.3690 ;
      RECT 0.0000 192.1490 37.2530 199.3690 ;
      RECT 0.0000 192.1490 38.1370 197.7710 ;
      RECT 0.0000 190.5490 37.2380 192.1490 ;
      RECT 0.0000 188.9530 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 183.3300 38.1370 188.9530 ;
      RECT 0.0000 181.7310 37.2400 183.3300 ;
      RECT 0.0000 180.1310 37.2370 181.7310 ;
      RECT 0.0000 30.2920 38.1370 180.1310 ;
      RECT 0.0000 28.6920 37.2370 30.2920 ;
      RECT 0.0000 18.2630 38.1370 28.6920 ;
      RECT 0.0000 16.1970 37.2370 18.2630 ;
      RECT 0.0000 10.7900 38.1370 16.1970 ;
      RECT 0.0000 9.1900 37.2370 10.7900 ;
      RECT 0.0000 0.9000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 0.9000 ;
      RECT 29.3550 246.8760 33.9550 246.8800 ;
      RECT 29.3550 0.0000 33.9550 246.8800 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1.2580 0.9000 ;
      RECT 36.6360 225.1960 38.1370 226.7820 ;
      RECT 0.0000 200.9690 38.1370 206.5930 ;
      RECT 0.0000 192.1490 37.2400 206.5930 ;
      RECT 0.0000 181.7310 37.2380 206.5930 ;
      RECT 0.0000 199.3690 37.2400 200.9690 ;
      RECT 0.0000 197.7710 37.2530 199.3690 ;
      RECT 0.0000 192.1490 37.2530 199.3690 ;
      RECT 0.0000 192.1490 38.1370 197.7710 ;
      RECT 0.0000 190.5490 37.2380 192.1490 ;
      RECT 0.0000 188.9530 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 183.3300 38.1370 188.9530 ;
      RECT 0.0000 181.7310 37.2400 183.3300 ;
      RECT 0.0000 180.1310 37.2370 181.7310 ;
      RECT 0.0000 30.2920 38.1370 180.1310 ;
      RECT 0.0000 28.6920 37.2370 30.2920 ;
      RECT 0.0000 18.2630 38.1370 28.6920 ;
      RECT 0.0000 16.1970 37.2370 18.2630 ;
      RECT 0.0000 10.7900 38.1370 16.1970 ;
      RECT 0.0000 9.1900 37.2370 10.7900 ;
      RECT 0.0000 0.9000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 0.9000 ;
      RECT 0.0000 228.3820 38.1370 247.8820 ;
      RECT 0.0000 208.1930 37.2430 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 223.2160 37.2430 228.3820 ;
      RECT 0.0000 208.1930 38.1370 223.2160 ;
      RECT 0.0000 206.5930 37.2370 208.1930 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1.2580 0.9000 ;
      RECT 36.6360 225.1960 38.1370 226.7820 ;
      RECT 0.0000 200.9690 38.1370 206.5930 ;
      RECT 0.0000 192.1490 37.2400 206.5930 ;
      RECT 0.0000 181.7310 37.2380 206.5930 ;
      RECT 0.0000 199.3690 37.2400 200.9690 ;
      RECT 0.0000 197.7710 37.2530 199.3690 ;
      RECT 0.0000 192.1490 37.2530 199.3690 ;
      RECT 0.0000 192.1490 38.1370 197.7710 ;
      RECT 0.0000 190.5490 37.2380 192.1490 ;
      RECT 0.0000 188.9530 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 181.7310 37.2400 190.5490 ;
      RECT 0.0000 183.3300 38.1370 188.9530 ;
      RECT 0.0000 181.7310 37.2400 183.3300 ;
      RECT 0.0000 180.1310 37.2370 181.7310 ;
      RECT 0.0000 30.2920 38.1370 180.1310 ;
      RECT 0.0000 28.6920 37.2370 30.2920 ;
      RECT 0.0000 18.2630 38.1370 28.6920 ;
      RECT 0.0000 16.1970 37.2370 18.2630 ;
      RECT 0.0000 10.7900 38.1370 16.1970 ;
      RECT 0.0000 9.1900 37.2370 10.7900 ;
      RECT 0.0000 0.9000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 9.1900 ;
      RECT 13.8010 0.0000 38.1370 0.9000 ;
      RECT 0.0000 228.3820 38.1370 247.8820 ;
      RECT 0.0000 208.1930 37.2430 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 0.9000 37.2370 247.8820 ;
      RECT 0.0000 223.2160 37.2430 228.3820 ;
      RECT 0.0000 208.1930 38.1370 223.2160 ;
      RECT 0.0000 206.5930 37.2370 208.1930 ;
  END
END SRAMLP1RW256x8

MACRO SRAMLP1RW256x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 110.509 BY 257.295 ;
  SYMMETRY X Y R90 ;

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.8580 0.0000 87.0580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.8580 0.0000 87.0580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.8580 0.0000 87.0580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.8580 0.0000 87.0580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.8580 0.0000 87.0580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.8970 0.0000 89.0970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.8970 0.0000 89.0970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.8970 0.0000 89.0970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.8970 0.0000 89.0970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.8970 0.0000 89.0970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[1]

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 42.1330 110.5090 42.3330 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 42.1330 110.5090 42.3330 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 42.1330 110.5090 42.3330 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 42.1330 110.5090 42.3330 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 42.1330 110.5090 42.3330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 3.1810 256.9950 3.4820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2800 256.9950 2.5790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.4800 256.9950 0.7800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3810 256.9950 1.6810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9800 256.9950 5.2800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.7800 256.9950 7.0790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8810 256.9950 6.1810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.6810 256.9950 7.9820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.0800 256.9950 4.3800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1810 256.9950 12.4800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.4800 256.9950 9.7800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.5800 256.9950 8.8800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.3810 256.9950 10.6810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.2810 256.9950 11.5810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.0810 256.9950 13.3800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.8800 256.9950 15.1810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.9800 256.9950 14.2810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.7800 256.9950 16.0800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.6800 256.9950 16.9800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.5810 256.9950 17.8810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.1800 256.9950 21.4800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.9800 256.9950 23.2790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.0810 256.9950 22.3810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.3810 256.9950 19.6820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.2800 256.9950 20.5800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4800 256.9950 18.7790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.6800 256.9950 25.9800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.7800 256.9950 25.0800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.8810 256.9950 24.1820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.5810 256.9950 26.8810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.4810 256.9950 27.7810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.0800 256.9950 31.3810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.3810 256.9950 28.6800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.1800 256.9950 30.4810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.9800 256.9950 32.2800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.2810 256.9950 29.5800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.3800 256.9950 37.6800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.5810 256.9950 35.8820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.4800 256.9950 36.7800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.6800 256.9950 34.9790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.8800 256.9950 33.1800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.7810 256.9950 34.0810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.1800 256.9950 39.4790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.2810 256.9950 38.5810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.8800 256.9950 42.1800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.9800 256.9950 41.2800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.0810 256.9950 40.3820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.5810 256.9950 44.8800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.3800 256.9950 46.6810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.7810 256.9950 43.0810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.6810 256.9950 43.9810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.4810 256.9950 45.7800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.2800 256.9950 47.5810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.7810 256.9950 52.0820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.1800 256.9950 48.4800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.8800 256.9950 51.1790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.0800 256.9950 49.3800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.9810 256.9950 50.2810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.5800 256.9950 53.8800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.3800 256.9950 55.6790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.4810 256.9950 54.7810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.2810 256.9950 56.5820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.6800 256.9950 52.9800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.7810 256.9950 61.0800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.0800 256.9950 58.3800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.1800 256.9950 57.4800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.9810 256.9950 59.2810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.8810 256.9950 60.1810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.4800 256.9950 63.7810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.5800 256.9950 62.8810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.3800 256.9950 64.6800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.6810 256.9950 61.9800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.2800 256.9950 65.5800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.1810 256.9950 66.4810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.7800 256.9950 70.0800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.6810 256.9950 70.9810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.9810 256.9950 68.2820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.8800 256.9950 69.1800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.0800 256.9950 67.3790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.5800 256.9950 71.8790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.2800 256.9950 74.5800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.3800 256.9950 73.6800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.4810 256.9950 72.7820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.1810 256.9950 75.4810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.6800 256.9950 79.9810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.9810 256.9950 77.2800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.7800 256.9950 79.0810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.5800 256.9950 80.8800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.0810 256.9950 76.3810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.8810 256.9950 78.1800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.1810 256.9950 84.4820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.0800 256.9950 85.3800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.2800 256.9950 83.5790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.4800 256.9950 81.7800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.3810 256.9950 82.6810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.9800 256.9950 86.2800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.7800 256.9950 88.0790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.8810 256.9950 87.1810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.5800 256.9950 89.8800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.6810 256.9950 88.9820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.1810 256.9950 93.4800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.4800 256.9950 90.7800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.9800 256.9950 95.2810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.3810 256.9950 91.6810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.2810 256.9950 92.5810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.0810 256.9950 94.3800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.8800 256.9950 96.1810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.7800 256.9950 97.0800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.4800 256.9950 99.7790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.6800 256.9950 97.9800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.5810 256.9950 98.8810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.1800 256.9950 102.4800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.9800 256.9950 104.2790 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.0810 256.9950 103.3810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.3810 256.9950 100.6820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.4810 256.9950 108.7810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.5810 256.9950 107.8810 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.8810 256.9950 105.1820 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.7800 256.9950 106.0800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.6800 256.9950 106.9800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.3810 256.9950 109.6800 257.2950 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.2800 256.9950 101.5800 257.2950 ;
    END
  END VSS

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 16.3970 110.5090 16.5970 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 16.3970 110.5090 16.5970 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 16.3970 110.5090 16.5970 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 16.3970 110.5090 16.5970 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 16.3970 110.5090 16.5970 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 16.8830 110.5090 17.0830 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 16.8830 110.5090 17.0830 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 16.8830 110.5090 17.0830 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 16.8830 110.5090 17.0830 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 16.8830 110.5090 17.0830 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 193.5870 110.5090 193.7870 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 193.5870 110.5090 193.7870 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 193.5870 110.5090 193.7870 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 193.5870 110.5090 193.7870 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 193.5870 110.5090 193.7870 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3150 239.5180 110.5090 239.7180 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3150 239.5180 110.5090 239.7180 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3150 239.5180 110.5090 239.7180 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3150 239.5180 110.5090 239.7180 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3150 239.5180 110.5090 239.7180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3150 235.9810 110.5090 236.1810 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3150 235.9810 110.5090 236.1810 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3150 235.9810 110.5090 236.1810 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3150 235.9810 110.5090 236.1810 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3150 235.9810 110.5090 236.1810 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3150 236.4740 110.5090 236.6740 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3150 236.4740 110.5090 236.6740 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3150 236.4740 110.5090 236.6740 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3150 236.4740 110.5090 236.6740 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3150 236.4740 110.5090 236.6740 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 96.3300 256.9920 96.6300 257.2920 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.2310 256.9920 97.5300 257.2920 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.1310 256.9920 98.4320 257.2920 ;
    END
    ANTENNADIFFAREA 7.0452 LAYER M5 ;
    ANTENNADIFFAREA 7.0452 LAYER M6 ;
    ANTENNADIFFAREA 7.0452 LAYER M7 ;
    ANTENNADIFFAREA 7.0452 LAYER M8 ;
    ANTENNADIFFAREA 7.0452 LAYER M9 ;
    ANTENNADIFFAREA 7.0452 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 230.8461 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 230.8461 LAYER M5 ;
  END VDDL

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.8180 0.0000 46.0180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.8180 0.0000 46.0180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.8180 0.0000 46.0180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.8180 0.0000 46.0180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.8180 0.0000 46.0180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.4850 0.0000 46.6850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.4850 0.0000 46.6850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.4850 0.0000 46.6850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.4850 0.0000 46.6850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.4850 0.0000 46.6850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[23]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.1860 0.0000 47.3860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.1860 0.0000 47.3860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.1860 0.0000 47.3860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.1860 0.0000 47.3860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.1860 0.0000 47.3860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.8530 0.0000 48.0530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.8530 0.0000 48.0530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.8530 0.0000 48.0530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.8530 0.0000 48.0530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.8530 0.0000 48.0530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[24]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.5540 0.0000 48.7540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.5540 0.0000 48.7540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.5540 0.0000 48.7540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.5540 0.0000 48.7540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.5540 0.0000 48.7540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.6020 0.0000 63.8020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.6020 0.0000 63.8020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.6020 0.0000 63.8020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.6020 0.0000 63.8020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.6020 0.0000 63.8020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.2340 0.0000 62.4340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.2340 0.0000 62.4340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.2340 0.0000 62.4340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.2340 0.0000 62.4340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.8660 0.0000 61.0660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.8660 0.0000 61.0660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.8660 0.0000 61.0660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.8660 0.0000 61.0660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.8660 0.0000 61.0660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.4980 0.0000 59.6980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.4980 0.0000 59.6980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.4980 0.0000 59.6980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.4980 0.0000 59.6980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.4980 0.0000 59.6980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.8040 0.0000 59.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.8040 0.0000 59.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.8040 0.0000 59.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.8040 0.0000 59.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.8040 0.0000 59.0040 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[19]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.4360 0.0000 57.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.4360 0.0000 57.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.4360 0.0000 57.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.4360 0.0000 57.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.4360 0.0000 57.6360 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[21]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.1300 0.0000 58.3300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.1300 0.0000 58.3300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.1300 0.0000 58.3300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.1300 0.0000 58.3300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.1300 0.0000 58.3300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.0620 0.0000 56.2620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.0620 0.0000 56.2620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.0620 0.0000 56.2620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.0620 0.0000 56.2620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.0620 0.0000 56.2620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[22]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.7620 0.0000 56.9620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.7620 0.0000 56.9620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.7620 0.0000 56.9620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.7620 0.0000 56.9620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.7620 0.0000 56.9620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.3940 0.0000 55.5940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.3940 0.0000 55.5940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.3940 0.0000 55.5940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.3940 0.0000 55.5940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.3940 0.0000 55.5940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.0260 0.0000 54.2260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.0260 0.0000 54.2260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.0260 0.0000 54.2260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.0260 0.0000 54.2260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.0260 0.0000 54.2260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.3250 0.0000 53.5250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.3250 0.0000 53.5250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.3250 0.0000 53.5250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.3250 0.0000 53.5250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.3250 0.0000 53.5250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[29]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.6970 0.0000 54.8970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.6970 0.0000 54.8970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.6970 0.0000 54.8970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.6970 0.0000 54.8970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.6970 0.0000 54.8970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[27]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.6580 0.0000 52.8580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.6580 0.0000 52.8580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.6580 0.0000 52.8580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.6580 0.0000 52.8580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.6580 0.0000 52.8580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.5890 0.0000 50.7890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.5890 0.0000 50.7890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.5890 0.0000 50.7890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.5890 0.0000 50.7890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.5890 0.0000 50.7890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[26]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.2900 0.0000 51.4900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.2900 0.0000 51.4900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.2900 0.0000 51.4900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.2900 0.0000 51.4900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.2900 0.0000 51.4900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.9220 0.0000 50.1220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.9220 0.0000 50.1220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.9220 0.0000 50.1220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.9220 0.0000 50.1220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.9220 0.0000 50.1220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.9570 0.0000 52.1570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.9570 0.0000 52.1570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.9570 0.0000 52.1570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.9570 0.0000 52.1570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.9570 0.0000 52.1570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M2 ;
  END O[28]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.2210 0.0000 49.4210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.2210 0.0000 49.4210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.2210 0.0000 49.4210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.2210 0.0000 49.4210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.2210 0.0000 49.4210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[25]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.8440 0.0000 74.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.8440 0.0000 74.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.8440 0.0000 74.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.8440 0.0000 74.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.8440 0.0000 74.0440 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[11]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.1780 0.0000 73.3780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.1780 0.0000 73.3780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.1780 0.0000 73.3780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.1780 0.0000 73.3780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.1780 0.0000 73.3780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.4800 0.0000 72.6800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.4800 0.0000 72.6800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.4800 0.0000 72.6800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.4800 0.0000 72.6800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.4800 0.0000 72.6800 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[8]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.1090 0.0000 71.3090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.1090 0.0000 71.3090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.1090 0.0000 71.3090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.1090 0.0000 71.3090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.1090 0.0000 71.3090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[7]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.5460 0.0000 74.7460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.5460 0.0000 74.7460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.5460 0.0000 74.7460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.5460 0.0000 74.7460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.5460 0.0000 74.7460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.4420 0.0000 70.6420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.4420 0.0000 70.6420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.4420 0.0000 70.6420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.4420 0.0000 70.6420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4420 0.0000 70.6420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.8100 0.0000 72.0100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.8100 0.0000 72.0100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.8100 0.0000 72.0100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.8100 0.0000 72.0100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.8100 0.0000 72.0100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.7410 0.0000 69.9410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.7410 0.0000 69.9410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.7410 0.0000 69.9410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.7410 0.0000 69.9410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.7410 0.0000 69.9410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[6]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.6370 0.0000 65.8370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.6370 0.0000 65.8370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.6370 0.0000 65.8370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.6370 0.0000 65.8370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6370 0.0000 65.8370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[4]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.3380 0.0000 66.5380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.3380 0.0000 66.5380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.3380 0.0000 66.5380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.3380 0.0000 66.5380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.3380 0.0000 66.5380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.9700 0.0000 65.1700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.9700 0.0000 65.1700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.9700 0.0000 65.1700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.9700 0.0000 65.1700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.9700 0.0000 65.1700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.0030 0.0000 67.2030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.0030 0.0000 67.2030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.0030 0.0000 67.2030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.0030 0.0000 67.2030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.0030 0.0000 67.2030 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[31]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.0740 0.0000 69.2740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.0740 0.0000 69.2740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.0740 0.0000 69.2740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.0740 0.0000 69.2740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.0740 0.0000 69.2740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.7060 0.0000 67.9060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.7060 0.0000 67.9060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.7060 0.0000 67.9060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.7060 0.0000 67.9060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.7060 0.0000 67.9060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3720 0.0000 68.5720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.3720 0.0000 68.5720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.3720 0.0000 68.5720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.3720 0.0000 68.5720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.3720 0.0000 68.5720 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[5]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.2670 0.0000 64.4670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.2670 0.0000 64.4670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.2670 0.0000 64.4670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.2670 0.0000 64.4670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.2670 0.0000 64.4670 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M2 ;
  END O[30]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.9010 0.0000 63.1010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.9010 0.0000 63.1010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.9010 0.0000 63.1010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.9010 0.0000 63.1010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.9010 0.0000 63.1010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[3]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.5330 0.0000 61.7330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.5330 0.0000 61.7330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.5330 0.0000 61.7330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.5330 0.0000 61.7330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.5330 0.0000 61.7330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[9]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.1650 0.0000 60.3650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.1650 0.0000 60.3650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.1650 0.0000 60.3650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.1650 0.0000 60.3650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.1650 0.0000 60.3650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[10]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 9.6830 110.5090 9.8830 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 9.6830 110.5090 9.8830 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 9.6830 110.5090 9.8830 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 9.6830 110.5090 9.8830 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 9.6830 110.5090 9.8830 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.1590 0.0000 86.3590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.1590 0.0000 86.3590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.1600 0.0000 86.3600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.1600 0.0000 86.3600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.1600 0.0000 86.3600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[2]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.7890 0.0000 84.9890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.7890 0.0000 84.9890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.7890 0.0000 84.9890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.7890 0.0000 84.9890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.7890 0.0000 84.9890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[20]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.4200 0.0000 83.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.4200 0.0000 83.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.4200 0.0000 83.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.4200 0.0000 83.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.4200 0.0000 83.6200 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[18]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.0520 0.0000 82.2520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.0520 0.0000 82.2520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.0520 0.0000 82.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.0520 0.0000 82.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.0520 0.0000 82.2520 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[17]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.4900 0.0000 85.6900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.4900 0.0000 85.6900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.4900 0.0000 85.6900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.4900 0.0000 85.6900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.4900 0.0000 85.6900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.1220 0.0000 84.3220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.1220 0.0000 84.3220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.1220 0.0000 84.3220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.1220 0.0000 84.3220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.1220 0.0000 84.3220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.7540 0.0000 82.9540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.7540 0.0000 82.9540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.7540 0.0000 82.9540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.7540 0.0000 82.9540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.7540 0.0000 82.9540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.3860 0.0000 81.5860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.3860 0.0000 81.5860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.3860 0.0000 81.5860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.3860 0.0000 81.5860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.3860 0.0000 81.5860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.6840 0.0000 80.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.6840 0.0000 80.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.6840 0.0000 80.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.6840 0.0000 80.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.6840 0.0000 80.8840 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[16]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.0180 0.0000 80.2180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.0180 0.0000 80.2180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.0180 0.0000 80.2180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.0180 0.0000 80.2180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.0180 0.0000 80.2180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.6500 0.0000 78.8500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.6500 0.0000 78.8500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.6500 0.0000 78.8500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.6500 0.0000 78.8500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.6500 0.0000 78.8500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.9140 0.0000 76.1140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.9140 0.0000 76.1140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.9140 0.0000 76.1140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.9140 0.0000 76.1140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.9140 0.0000 76.1140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.2820 0.0000 77.4820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.2820 0.0000 77.4820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.2820 0.0000 77.4820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.2820 0.0000 77.4820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.2820 0.0000 77.4820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.3170 0.0000 79.5170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.3170 0.0000 79.5170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.3170 0.0000 79.5170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.3170 0.0000 79.5170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.3170 0.0000 79.5170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[15]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.9510 0.0000 78.1510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.9510 0.0000 78.1510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.9510 0.0000 78.1510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.9510 0.0000 78.1510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.9510 0.0000 78.1510 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[14]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.5830 0.0000 76.7830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.5830 0.0000 76.7830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.5830 0.0000 76.7830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.5830 0.0000 76.7830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.5830 0.0000 76.7830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1538 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1538 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1538 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1538 LAYER M2 ;
  END O[13]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.2120 0.0000 75.4120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.2120 0.0000 75.4120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.2120 0.0000 75.4120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.2120 0.0000 75.4120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2120 0.0000 75.4120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[12]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 220.0470 110.5090 220.2470 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 220.0470 110.5090 220.2470 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 220.0470 110.5090 220.2470 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 220.0470 110.5090 220.2470 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 220.0470 110.5090 220.2470 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.5820 0.0000 89.7820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.5820 0.0000 89.7820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.5820 0.0000 89.7820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.5820 0.0000 89.7820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.5820 0.0000 89.7820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 211.2270 110.5090 211.4270 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 211.2270 110.5090 211.4270 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 211.2270 110.5090 211.4270 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 211.2270 110.5090 211.4270 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 211.2270 110.5090 211.4270 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 212.8170 110.5090 213.0170 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 212.8170 110.5090 213.0170 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 212.8170 110.5090 213.0170 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 212.8170 110.5090 213.0170 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 212.8170 110.5090 213.0170 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 104.4300 256.9920 104.7300 257.2920 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.2300 256.9920 106.5290 257.2920 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.3310 256.9920 105.6310 257.2920 ;
    END
  END VDD

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 203.9970 110.5090 204.1970 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 203.9970 110.5090 204.1970 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 203.9970 110.5090 204.1970 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 203.9970 110.5090 204.1970 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 203.9970 110.5090 204.1970 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 202.4070 110.5090 202.6070 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 202.4070 110.5090 202.6070 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 202.4070 110.5090 202.6070 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 202.4070 110.5090 202.6070 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 202.4070 110.5090 202.6070 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3090 195.1770 110.5090 195.3770 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3090 195.1770 110.5090 195.3770 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3090 195.1770 110.5090 195.3770 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3090 195.1770 110.5090 195.3770 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3090 195.1770 110.5090 195.3770 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.2260 0.0000 88.4260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.2260 0.0000 88.4260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.2260 0.0000 88.4260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.2260 0.0000 88.4260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.2260 0.0000 88.4260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.5230 0.0000 87.7230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.5230 0.0000 87.7230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.5230 0.0000 87.7230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.5230 0.0000 87.7230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.5230 0.0000 87.7230 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[0]
  OBS
    LAYER M2 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 235.2810 109.6150 240.4180 ;
      RECT 0.0000 220.9470 110.5090 235.2810 ;
      RECT 0.0000 219.3470 109.6090 220.9470 ;
      RECT 109.6150 237.3740 110.5090 238.8180 ;
      RECT 0.0000 213.7170 110.5090 219.3470 ;
      RECT 0.0000 210.5270 109.6090 213.7170 ;
      RECT 0.0000 204.8970 110.5090 210.5270 ;
      RECT 0.0000 201.7070 109.6090 204.8970 ;
      RECT 0.0000 196.0770 110.5090 201.7070 ;
      RECT 0.0000 192.8870 109.6090 196.0770 ;
      RECT 0.0000 43.0330 110.5090 192.8870 ;
      RECT 0.0000 41.4330 109.6090 43.0330 ;
      RECT 0.0000 17.7830 110.5090 41.4330 ;
      RECT 0.0000 15.6970 109.6090 17.7830 ;
      RECT 0.0000 10.5830 110.5090 15.6970 ;
      RECT 0.0000 8.9830 109.6090 10.5830 ;
      RECT 0.0000 0.9000 110.5090 8.9830 ;
      RECT 0.0000 0.0000 45.1180 0.9000 ;
      RECT 90.4820 0.0000 110.5090 8.9830 ;
      RECT 90.4820 0.0000 110.5090 0.9000 ;
      RECT 0.0000 240.4180 110.5090 257.2950 ;
      RECT 0.0000 220.9470 109.6150 257.2950 ;
      RECT 0.0000 0.0000 45.1180 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
    LAYER M1 ;
      RECT 109.7090 212.0270 110.5090 212.2170 ;
      RECT 109.7090 203.2070 110.5090 203.3970 ;
      RECT 109.7090 194.3870 110.5090 194.5770 ;
      RECT 109.0080 237.2740 110.5090 238.9180 ;
      RECT 0.0000 213.6170 110.5090 219.4470 ;
      RECT 0.0000 210.6270 109.7090 213.6170 ;
      RECT 0.0000 204.7970 110.5090 210.6270 ;
      RECT 0.0000 201.8070 109.7090 204.7970 ;
      RECT 0.0000 195.9770 110.5090 201.8070 ;
      RECT 0.0000 192.9870 109.7090 195.9770 ;
      RECT 0.0000 42.9330 110.5090 192.9870 ;
      RECT 0.0000 41.5330 109.7090 42.9330 ;
      RECT 0.0000 17.6830 110.5090 41.5330 ;
      RECT 0.0000 15.7970 109.7090 17.6830 ;
      RECT 0.0000 10.4830 110.5090 15.7970 ;
      RECT 0.0000 9.0830 109.7090 10.4830 ;
      RECT 0.0000 0.8000 110.5090 9.0830 ;
      RECT 0.0000 0.0000 45.2180 0.8000 ;
      RECT 90.3820 0.0000 110.5090 9.0830 ;
      RECT 90.3820 0.0000 110.5090 0.8000 ;
      RECT 0.0000 240.3180 110.5090 257.2950 ;
      RECT 0.0000 220.8470 109.7150 257.2950 ;
      RECT 0.0000 0.0000 45.2180 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 0.8000 109.7090 257.2950 ;
      RECT 0.0000 235.3810 109.7150 240.3180 ;
      RECT 0.0000 220.8470 110.5090 235.3810 ;
      RECT 0.0000 219.4470 109.7090 220.8470 ;
    LAYER PO ;
      RECT 0.0000 0.0000 110.5090 257.2950 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 110.5090 257.2950 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 110.5090 257.2950 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 110.5090 257.2950 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 110.5090 257.2950 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 110.5090 257.2950 ;
    LAYER M5 ;
      RECT 110.3800 256.2950 110.5090 257.2950 ;
      RECT 109.6150 237.3740 110.5090 238.8180 ;
      RECT 107.2290 256.2920 110.5090 256.2950 ;
      RECT 107.2290 240.4180 110.5090 256.2950 ;
      RECT 99.1320 256.2920 103.7300 256.2950 ;
      RECT 99.1320 0.0000 103.7300 256.2950 ;
      RECT 0.0000 256.2920 95.6300 256.2950 ;
      RECT 0.0000 0.9000 95.6300 256.2950 ;
      RECT 0.0000 0.0000 45.1180 256.2920 ;
      RECT 0.0000 240.4180 110.5090 256.2920 ;
      RECT 0.0000 220.9470 109.6150 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 0.9000 109.6090 256.2920 ;
      RECT 0.0000 235.2810 109.6150 240.4180 ;
      RECT 0.0000 220.9470 110.5090 235.2810 ;
      RECT 0.0000 219.3470 109.6090 220.9470 ;
      RECT 0.0000 213.7170 110.5090 219.3470 ;
      RECT 0.0000 210.5270 109.6090 213.7170 ;
      RECT 0.0000 204.8970 110.5090 210.5270 ;
      RECT 0.0000 201.7070 109.6090 204.8970 ;
      RECT 0.0000 196.0770 110.5090 201.7070 ;
      RECT 0.0000 192.8870 109.6090 196.0770 ;
      RECT 0.0000 43.0330 110.5090 192.8870 ;
      RECT 0.0000 41.4330 109.6090 43.0330 ;
      RECT 0.0000 17.7830 110.5090 41.4330 ;
      RECT 0.0000 15.6970 109.6090 17.7830 ;
      RECT 0.0000 10.5830 110.5090 15.6970 ;
      RECT 0.0000 8.9830 109.6090 10.5830 ;
      RECT 0.0000 0.9000 110.5090 8.9830 ;
      RECT 0.0000 0.0000 45.1180 0.9000 ;
      RECT 90.4820 0.0000 110.5090 8.9830 ;
      RECT 90.4820 0.0000 110.5090 0.9000 ;
    LAYER M4 ;
      RECT 109.6150 237.3740 110.5090 238.8180 ;
      RECT 0.0000 213.7170 110.5090 219.3470 ;
      RECT 0.0000 210.5270 109.6090 213.7170 ;
      RECT 0.0000 204.8970 110.5090 210.5270 ;
      RECT 0.0000 201.7070 109.6090 204.8970 ;
      RECT 0.0000 196.0770 110.5090 201.7070 ;
      RECT 0.0000 192.8870 109.6090 196.0770 ;
      RECT 0.0000 43.0330 110.5090 192.8870 ;
      RECT 0.0000 41.4330 109.6090 43.0330 ;
      RECT 0.0000 17.7830 110.5090 41.4330 ;
      RECT 0.0000 15.6970 109.6090 17.7830 ;
      RECT 0.0000 10.5830 110.5090 15.6970 ;
      RECT 0.0000 8.9830 109.6090 10.5830 ;
      RECT 0.0000 0.9000 110.5090 8.9830 ;
      RECT 0.0000 0.0000 45.1180 0.9000 ;
      RECT 90.4820 0.0000 110.5090 8.9830 ;
      RECT 90.4820 0.0000 110.5090 0.9000 ;
      RECT 0.0000 240.4180 110.5090 257.2950 ;
      RECT 0.0000 220.9470 109.6150 257.2950 ;
      RECT 0.0000 0.0000 45.1180 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 235.2810 109.6150 240.4180 ;
      RECT 0.0000 220.9470 110.5090 235.2810 ;
      RECT 0.0000 219.3470 109.6090 220.9470 ;
    LAYER M3 ;
      RECT 109.6150 237.3740 110.5090 238.8180 ;
      RECT 0.0000 213.7170 110.5090 219.3470 ;
      RECT 0.0000 210.5270 109.6090 213.7170 ;
      RECT 0.0000 204.8970 110.5090 210.5270 ;
      RECT 0.0000 201.7070 109.6090 204.8970 ;
      RECT 0.0000 196.0770 110.5090 201.7070 ;
      RECT 0.0000 192.8870 109.6090 196.0770 ;
      RECT 0.0000 43.0330 110.5090 192.8870 ;
      RECT 0.0000 41.4330 109.6090 43.0330 ;
      RECT 0.0000 17.7830 110.5090 41.4330 ;
      RECT 0.0000 15.6970 109.6090 17.7830 ;
      RECT 0.0000 10.5830 110.5090 15.6970 ;
      RECT 0.0000 8.9830 109.6090 10.5830 ;
      RECT 0.0000 0.9000 110.5090 8.9830 ;
      RECT 0.0000 0.0000 45.1180 0.9000 ;
      RECT 90.4820 0.0000 110.5090 8.9830 ;
      RECT 90.4820 0.0000 110.5090 0.9000 ;
      RECT 0.0000 240.4180 110.5090 257.2950 ;
      RECT 0.0000 220.9470 109.6150 257.2950 ;
      RECT 0.0000 0.0000 45.1180 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 0.9000 109.6090 257.2950 ;
      RECT 0.0000 235.2810 109.6150 240.4180 ;
      RECT 0.0000 220.9470 110.5090 235.2810 ;
      RECT 0.0000 219.3470 109.6090 220.9470 ;
  END
END SRAMLP1RW256x32

MACRO SRAMLP1RW256x46
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 148.491 BY 264.758 ;
  SYMMETRY X Y R90 ;

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.2880 0.0000 120.4880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.2880 0.0000 120.4880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.2880 0.0000 120.4880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.2880 0.0000 120.4880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.2880 0.0000 120.4880 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[16]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.5070 0.0000 89.7070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.5070 0.0000 89.7070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.5070 0.0000 89.7070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.5070 0.0000 89.7070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.5070 0.0000 89.7070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.8190 0.0000 102.0190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.8190 0.0000 102.0190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.8190 0.0000 102.0190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.8190 0.0000 102.0190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.8190 0.0000 102.0190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.1360 0.0000 101.3360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.1360 0.0000 101.3360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.1360 0.0000 101.3360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.1360 0.0000 101.3360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.1360 0.0000 101.3360 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[39]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.5550 0.0000 104.7550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.5550 0.0000 104.7550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.5550 0.0000 104.7550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.5550 0.0000 104.7550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.5550 0.0000 104.7550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8720 0.0000 104.0720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8720 0.0000 104.0720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8720 0.0000 104.0720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8720 0.0000 104.0720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8720 0.0000 104.0720 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[18]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6110 0.0000 93.8110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6110 0.0000 93.8110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6110 0.0000 93.8110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6110 0.0000 93.8110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6110 0.0000 93.8110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2970 243.5910 148.4910 243.7910 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2970 243.5910 148.4910 243.7910 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2970 243.5910 148.4910 243.7910 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2970 243.5910 148.4910 243.7910 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2970 243.5910 148.4910 243.7910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2970 246.9670 148.4910 247.1670 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2970 246.9670 148.4910 247.1670 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2970 246.9670 148.4910 247.1670 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2970 246.9670 148.4910 247.1670 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2970 246.9670 148.4910 247.1670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2940 220.5200 148.4910 220.7200 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2940 220.5200 148.4910 220.7200 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2940 220.5200 148.4910 220.7200 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2940 220.5200 148.4910 220.7200 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2940 220.5200 148.4910 220.7200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2910 227.7500 148.4910 227.9500 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2910 227.7500 148.4910 227.9500 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2910 227.7500 148.4910 227.9500 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2910 227.7500 148.4910 227.9500 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2910 227.7500 148.4910 227.9500 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.3070 218.9300 148.4910 219.1300 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.3070 218.9300 148.4910 219.1300 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.3070 218.9300 148.4910 219.1300 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.3070 218.9300 148.4910 219.1300 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.3070 218.9300 148.4910 219.1300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.0880 0.0000 86.2880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.0880 0.0000 86.2880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.0880 0.0000 86.2880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.0880 0.0000 86.2880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.0880 0.0000 86.2880 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[26]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.2910 0.0000 107.4910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.2910 0.0000 107.4910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.2910 0.0000 107.4910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.2910 0.0000 107.4910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.2910 0.0000 107.4910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.6080 0.0000 106.8080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.6080 0.0000 106.8080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.6080 0.0000 106.8080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.6080 0.0000 106.8080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.6080 0.0000 106.8080 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[41]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.7710 0.0000 86.9710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.7710 0.0000 86.9710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.7710 0.0000 86.9710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.7710 0.0000 86.9710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.7710 0.0000 86.9710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.9310 0.0000 80.1310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.9310 0.0000 80.1310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.9310 0.0000 80.1310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.9310 0.0000 80.1310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.9310 0.0000 80.1310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.2480 0.0000 79.4480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.2480 0.0000 79.4480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.2480 0.0000 79.4480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.2480 0.0000 79.4480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.2480 0.0000 79.4480 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[32]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.2990 0.0000 81.4990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.2990 0.0000 81.4990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.2990 0.0000 81.4990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.2990 0.0000 81.4990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.2990 0.0000 81.4990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2910 49.8360 148.4910 50.0360 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2910 49.8360 148.4910 50.0360 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2910 49.8360 148.4910 50.0360 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2910 49.8360 148.4910 50.0360 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2910 49.8360 148.4910 50.0360 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2910 9.8180 148.4910 10.0180 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2910 9.8180 148.4910 10.0180 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2910 9.8180 148.4910 10.0180 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2910 9.8180 148.4910 10.0180 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2910 9.8180 148.4910 10.0180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2910 17.2900 148.4910 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2910 17.2900 148.4910 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2910 17.2900 148.4910 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2910 17.2900 148.4910 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2910 17.2900 148.4910 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 139.0500 264.4580 139.3500 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.9490 264.4580 140.2480 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.8500 264.4580 141.1510 264.7580 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.8830 0.0000 65.0830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.8830 0.0000 65.0830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.8830 0.0000 65.0830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.8830 0.0000 65.0830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.8830 0.0000 65.0830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.3950 0.0000 111.5950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.3950 0.0000 111.5950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.3950 0.0000 111.5950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.3950 0.0000 111.5950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.3950 0.0000 111.5950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2940 202.8800 148.4910 203.0800 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2940 202.8800 148.4910 203.0800 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2940 202.8800 148.4910 203.0800 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2940 202.8800 148.4910 203.0800 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2940 202.8800 148.4910 203.0800 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2920 211.7000 148.4910 211.9000 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2920 211.7000 148.4910 211.9000 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2920 211.7000 148.4910 211.9000 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2920 211.7000 148.4910 211.9000 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2920 211.7000 148.4910 211.9000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2940 210.1100 148.4910 210.3100 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2940 210.1100 148.4910 210.3100 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2940 210.1100 148.4910 210.3100 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2940 210.1100 148.4910 210.3100 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2940 210.1100 148.4910 210.3100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2910 201.2900 148.4910 201.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2910 201.2900 148.4910 201.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2910 201.2900 148.4910 201.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2910 201.2900 148.4910 201.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2910 201.2900 148.4910 201.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2970 244.2150 148.4910 244.4150 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2970 244.2150 148.4910 244.4150 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2970 244.2150 148.4910 244.4150 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2970 244.2150 148.4910 244.4150 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2970 244.2150 148.4910 244.4150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 146.2490 264.4570 146.5490 264.7570 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.3500 264.4570 145.6510 264.7570 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.1490 264.4570 147.4500 264.7570 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 1.8000 264.4580 2.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.9000 264.4580 1.2000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 264.4580 0.3000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.3990 264.4580 5.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.5990 264.4580 3.9000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7000 264.4580 2.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.2000 264.4580 7.5000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.4990 264.4580 4.8000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.2990 264.4580 6.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.7990 264.4580 11.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7000 264.4580 12.0000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.0990 264.4580 8.3980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.8990 264.4580 10.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.0000 264.4580 9.3010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.2000 264.4580 16.5000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.3990 264.4580 14.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.5000 264.4580 13.8010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.5990 264.4580 12.8980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.2990 264.4580 15.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0000 264.4580 18.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1000 264.4580 17.4000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.5990 264.4580 21.8990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.7990 264.4580 20.1000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.9000 264.4580 19.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.6990 264.4580 21.0000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.4000 264.4580 23.7000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.2990 264.4580 24.5980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.0990 264.4580 26.3990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.2000 264.4580 25.5010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.4990 264.4580 22.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.9990 264.4580 27.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.5990 264.4580 30.8990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.9000 264.4580 28.2000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.7000 264.4580 30.0010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.7990 264.4580 29.0980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.2000 264.4580 34.4990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.3000 264.4580 33.6000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.9990 264.4580 36.3000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.4000 264.4580 32.7000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.1000 264.4580 35.3990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.4990 264.4580 31.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.7990 264.4580 38.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.6000 264.4580 39.9000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.4990 264.4580 40.7980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.8990 264.4580 37.2000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.6990 264.4580 38.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.1990 264.4580 43.4990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.1000 264.4580 44.4000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.9990 264.4580 45.2980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.2990 264.4580 42.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.4000 264.4580 41.7010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.4000 264.4580 50.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.5000 264.4580 49.8000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.7990 264.4580 47.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.9000 264.4580 46.2010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.6990 264.4580 47.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.6000 264.4580 48.9000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.9990 264.4580 54.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.1990 264.4580 52.5000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.3000 264.4580 51.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.0990 264.4580 53.4000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.8990 264.4580 55.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.3990 264.4580 59.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.8000 264.4580 56.1000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.3000 264.4580 60.6000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.6990 264.4580 56.9980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.4990 264.4580 58.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.6000 264.4580 57.9010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.9990 264.4580 63.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.1000 264.4580 62.4010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.1990 264.4580 61.4980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.8990 264.4580 64.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.8000 264.4580 65.1000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.6000 264.4580 66.8990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.7000 264.4580 66.0000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.3990 264.4580 68.7000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.5000 264.4580 67.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.2990 264.4580 69.6000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.1990 264.4580 70.4990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.0000 264.4580 72.3000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.8990 264.4580 73.1980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.6990 264.4580 74.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.8000 264.4580 74.1010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.0990 264.4580 71.3990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.5990 264.4580 75.8990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.1990 264.4580 79.4990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.5000 264.4580 76.8000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.3000 264.4580 78.6010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.3990 264.4580 77.6980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.8000 264.4580 83.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.9000 264.4580 82.2000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.7000 264.4580 83.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.0990 264.4580 80.3990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.0000 264.4580 81.3000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.3990 264.4580 86.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.5990 264.4580 84.9000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.2000 264.4580 88.5000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.0990 264.4580 89.3980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.4990 264.4580 85.8000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.2990 264.4580 87.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.7990 264.4580 92.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.7000 264.4580 93.0000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.5990 264.4580 93.8980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.8990 264.4580 91.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.0000 264.4580 90.3010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.1000 264.4580 98.4000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.3990 264.4580 95.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.5000 264.4580 94.8010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.2990 264.4580 96.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.2000 264.4580 97.5000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.0000 264.4580 99.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.5990 264.4580 102.8990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.7990 264.4580 101.1000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.9000 264.4580 100.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.6990 264.4580 102.0000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.4990 264.4580 103.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.9990 264.4580 108.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.4000 264.4580 104.7000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.2990 264.4580 105.5980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.0990 264.4580 107.3990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.2000 264.4580 106.5010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.5990 264.4580 111.8990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.9000 264.4580 109.2000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.7000 264.4580 111.0010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.7990 264.4580 110.0980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.4990 264.4580 112.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.2000 264.4580 115.4990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.3000 264.4580 114.6000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.9990 264.4580 117.3000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.1000 264.4580 116.3990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.8990 264.4580 118.2000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.4000 264.4580 113.7000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.7990 264.4580 119.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.6000 264.4580 120.9000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.4990 264.4580 121.7980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.4000 264.4580 122.7010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.6990 264.4580 119.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.1990 264.4580 124.4990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.1000 264.4580 125.4000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.9000 264.4580 127.2010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.9990 264.4580 126.2980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.2990 264.4580 123.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.5000 264.4580 130.8000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.3000 264.4580 132.5990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.7990 264.4580 128.0990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.4000 264.4580 131.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.6990 264.4580 128.9990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.6000 264.4580 129.9000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.9990 264.4580 135.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.1990 264.4580 133.5000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.8000 264.4580 137.1000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.0990 264.4580 134.4000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.8990 264.4580 136.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.3990 264.4580 140.6990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.3000 264.4580 141.6000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.6990 264.4580 137.9980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.4990 264.4580 139.7990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.8000 264.4580 146.1000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.8990 264.4580 145.1990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.1990 264.4580 142.4980 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.1000 264.4580 143.4010 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.9990 264.4580 144.2990 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.7000 264.4580 147.0000 264.7580 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.6000 264.4580 138.9010 264.7580 ;
    END
  END VSS

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 127.1280 0.0000 127.3280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.1280 0.0000 127.3280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.1280 0.0000 127.3280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 127.1280 0.0000 127.3280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 127.1280 0.0000 127.3280 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[7]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.6190 0.0000 67.8190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.6190 0.0000 67.8190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.6190 0.0000 67.8190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.6190 0.0000 67.8190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.6190 0.0000 67.8190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.9360 0.0000 67.1360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.9360 0.0000 67.1360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.9360 0.0000 67.1360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.9360 0.0000 67.1360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.9360 0.0000 67.1360 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[30]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4560 0.0000 87.6560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4560 0.0000 87.6560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4560 0.0000 87.6560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4560 0.0000 87.6560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4560 0.0000 87.6560 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[35]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 127.8000 0.0000 128.0000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.8000 0.0000 128.0000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.8000 0.0000 128.0000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 127.8000 0.0000 128.0000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 127.8000 0.0000 128.0000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.7230 0.0000 71.9230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.7230 0.0000 71.9230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.7230 0.0000 71.9230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.7230 0.0000 71.9230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.7230 0.0000 71.9230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.0400 0.0000 71.2400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.0400 0.0000 71.2400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.0400 0.0000 71.2400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.0400 0.0000 71.2400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.0400 0.0000 71.2400 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[34]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.9870 0.0000 69.1870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.9870 0.0000 69.1870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.9870 0.0000 69.1870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.9870 0.0000 69.1870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.9870 0.0000 69.1870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.2910 16.8280 148.4910 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.2910 16.8280 148.4910 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.2910 16.8280 148.4910 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.2910 16.8280 148.4910 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.2910 16.8280 148.4910 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7120 0.0000 110.9120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7120 0.0000 110.9120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7120 0.0000 110.9120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7120 0.0000 110.9120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7120 0.0000 110.9120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[11]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3040 0.0000 68.5040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.3040 0.0000 68.5040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.3040 0.0000 68.5040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.3040 0.0000 68.5040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.3040 0.0000 68.5040 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[2]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.7200 0.0000 84.9200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.7200 0.0000 84.9200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.7200 0.0000 84.9200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.7200 0.0000 84.9200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.7200 0.0000 84.9200 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[40]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.3520 0.0000 83.5520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.3520 0.0000 83.5520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.3520 0.0000 83.5520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.3520 0.0000 83.5520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.3520 0.0000 83.5520 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[27]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.4030 0.0000 85.6030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.4030 0.0000 85.6030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.4030 0.0000 85.6030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.4030 0.0000 85.6030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.4030 0.0000 85.6030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.9230 0.0000 106.1230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.9230 0.0000 106.1230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.9230 0.0000 106.1230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.9230 0.0000 106.1230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.9230 0.0000 106.1230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[41]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 113.4480 0.0000 113.6480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.4480 0.0000 113.6480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.4480 0.0000 113.6480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 113.4480 0.0000 113.6480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.4480 0.0000 113.6480 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[33]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.8670 0.0000 117.0670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.8670 0.0000 117.0670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.8670 0.0000 117.0670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.8670 0.0000 117.0670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.8670 0.0000 117.0670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 115.4990 0.0000 115.6990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.4990 0.0000 115.6990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.4990 0.0000 115.6990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.4990 0.0000 115.6990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.4990 0.0000 115.6990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.1840 0.0000 116.3840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.1840 0.0000 116.3840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.1840 0.0000 116.3840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.1840 0.0000 116.3840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.1840 0.0000 116.3840 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[9]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 118.9200 0.0000 119.1200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.9200 0.0000 119.1200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.9200 0.0000 119.1200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 118.9200 0.0000 119.1200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.9200 0.0000 119.1200 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[1]

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 114.8160 0.0000 115.0160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.8160 0.0000 115.0160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.8160 0.0000 115.0160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.8160 0.0000 115.0160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.8160 0.0000 115.0160 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[44]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 114.1310 0.0000 114.3310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.1310 0.0000 114.3310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.1310 0.0000 114.3310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.1310 0.0000 114.3310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.1310 0.0000 114.3310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 121.6560 0.0000 121.8560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.6560 0.0000 121.8560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.6560 0.0000 121.8560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 121.6560 0.0000 121.8560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.6560 0.0000 121.8560 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[3]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 122.3390 0.0000 122.5390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.3390 0.0000 122.5390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.3390 0.0000 122.5390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 122.3390 0.0000 122.5390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.3390 0.0000 122.5390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[42]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 124.3920 0.0000 124.5920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.3920 0.0000 124.5920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.3920 0.0000 124.5920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 124.3920 0.0000 124.5920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.3920 0.0000 124.5920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[4]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 125.0750 0.0000 125.2750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.0750 0.0000 125.2750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.0750 0.0000 125.2750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 125.0750 0.0000 125.2750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 125.0750 0.0000 125.2750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[37]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 119.6030 0.0000 119.8030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.6030 0.0000 119.8030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.6030 0.0000 119.8030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.6030 0.0000 119.8030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.6030 0.0000 119.8030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 125.7600 0.0000 125.9600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.7600 0.0000 125.9600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.7600 0.0000 125.9600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 125.7600 0.0000 125.9600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 125.7600 0.0000 125.9600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[37]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 126.4430 0.0000 126.6430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.4430 0.0000 126.6430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.4430 0.0000 126.6430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 126.4430 0.0000 126.6430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 126.4430 0.0000 126.6430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.7150 0.0000 97.9150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.7150 0.0000 97.9150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.7150 0.0000 97.9150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.7150 0.0000 97.9150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.7150 0.0000 97.9150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.5120 0.0000 76.7120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.5120 0.0000 76.7120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.5120 0.0000 76.7120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.5120 0.0000 76.7120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.5120 0.0000 76.7120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[5]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.0320 0.0000 97.2320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.0320 0.0000 97.2320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.0320 0.0000 97.2320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.0320 0.0000 97.2320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.0320 0.0000 97.2320 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[24]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.1950 0.0000 77.3950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.1950 0.0000 77.3950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.1950 0.0000 77.3950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.1950 0.0000 77.3950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.1950 0.0000 77.3950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.8800 0.0000 78.0800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.8800 0.0000 78.0800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.8800 0.0000 78.0800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.8800 0.0000 78.0800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.8800 0.0000 78.0800 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[15]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.3470 0.0000 96.5470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.3470 0.0000 96.5470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.3470 0.0000 96.5470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.3470 0.0000 96.5470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.3470 0.0000 96.5470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.6640 0.0000 95.8640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.6640 0.0000 95.8640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.6640 0.0000 95.8640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.6640 0.0000 95.8640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.6640 0.0000 95.8640 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[38]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.5630 0.0000 78.7630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.5630 0.0000 78.7630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.5630 0.0000 78.7630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.5630 0.0000 78.7630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.5630 0.0000 78.7630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.0830 0.0000 99.2830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.0830 0.0000 99.2830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.0830 0.0000 99.2830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.0830 0.0000 99.2830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.0830 0.0000 99.2830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.9790 0.0000 95.1790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.9790 0.0000 95.1790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.9790 0.0000 95.1790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.9790 0.0000 95.1790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.9790 0.0000 95.1790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.4000 0.0000 98.6000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.4000 0.0000 98.6000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.4000 0.0000 98.6000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.4000 0.0000 98.6000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.4000 0.0000 98.6000 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[31]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.7680 0.0000 99.9680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.7680 0.0000 99.9680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.7680 0.0000 99.9680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.7680 0.0000 99.9680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.7680 0.0000 99.9680 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[23]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.4510 0.0000 100.6510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.4510 0.0000 100.6510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.4510 0.0000 100.6510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.4510 0.0000 100.6510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.4510 0.0000 100.6510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[39]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.2960 0.0000 94.4960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.2960 0.0000 94.4960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.2960 0.0000 94.4960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.2960 0.0000 94.4960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.2960 0.0000 94.4960 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[13]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.8750 0.0000 91.0750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.8750 0.0000 91.0750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.8750 0.0000 91.0750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.8750 0.0000 91.0750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.8750 0.0000 91.0750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.2400 0.0000 105.4400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.2400 0.0000 105.4400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.2400 0.0000 105.4400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.2400 0.0000 105.4400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.2400 0.0000 105.4400 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[21]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.1920 0.0000 90.3920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.1920 0.0000 90.3920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.1920 0.0000 90.3920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.1920 0.0000 90.3920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.1920 0.0000 90.3920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[17]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.1390 0.0000 88.3390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.1390 0.0000 88.3390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.1390 0.0000 88.3390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.1390 0.0000 88.3390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.1390 0.0000 88.3390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.0350 0.0000 84.2350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.0350 0.0000 84.2350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.0350 0.0000 84.2350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.0350 0.0000 84.2350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.0350 0.0000 84.2350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[40]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.9280 0.0000 93.1280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.9280 0.0000 93.1280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.9280 0.0000 93.1280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.9280 0.0000 93.1280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.9280 0.0000 93.1280 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[36]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 112.7630 0.0000 112.9630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.7630 0.0000 112.9630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.7630 0.0000 112.9630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 112.7630 0.0000 112.9630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.7630 0.0000 112.9630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 112.0800 0.0000 112.2800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.0800 0.0000 112.2800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.0800 0.0000 112.2800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 112.0800 0.0000 112.2800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.0800 0.0000 112.2800 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[20]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.2510 0.0010 66.4510 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.2510 0.0010 66.4510 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.2510 0.0000 66.4510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.2510 0.0000 66.4510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.2510 0.0000 66.4510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.6590 0.0000 108.8590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.6590 0.0000 108.8590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.6590 0.0000 108.8590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.6590 0.0000 108.8590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.6590 0.0000 108.8590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5680 0.0000 65.7680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5680 0.0000 65.7680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5680 0.0000 65.7680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5680 0.0000 65.7680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5680 0.0000 65.7680 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[0]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.6720 0.0000 69.8720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.6720 0.0000 69.8720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.6720 0.0000 69.8720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.6720 0.0000 69.8720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.6720 0.0000 69.8720 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[19]

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.3440 0.0000 109.5440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.3440 0.0000 109.5440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.3440 0.0000 109.5440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.3440 0.0000 109.5440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.3440 0.0000 109.5440 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[45]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.0270 0.0000 110.2270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.0270 0.0000 110.2270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.0270 0.0000 110.2270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.0270 0.0000 110.2270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.0270 0.0000 110.2270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.3550 0.0000 70.5550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.3550 0.0000 70.5550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.3550 0.0000 70.5550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.3550 0.0000 70.5550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.3550 0.0000 70.5550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.9760 0.0000 108.1760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.9760 0.0000 108.1760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.9760 0.0000 108.1760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.9760 0.0000 108.1760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.9760 0.0000 108.1760 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[12]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.0910 0.0000 73.2910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.0910 0.0000 73.2910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.0910 0.0000 73.2910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.0910 0.0000 73.2910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.0910 0.0000 73.2910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.4080 0.0000 72.6080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.4080 0.0000 72.6080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.4080 0.0000 72.6080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.4080 0.0000 72.6080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.4080 0.0000 72.6080 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[29]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.7760 0.0000 73.9760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.7760 0.0000 73.9760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.7760 0.0000 73.9760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.7760 0.0000 73.9760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.7760 0.0000 73.9760 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[43]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.1870 0.0000 103.3870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.1870 0.0000 103.3870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.1870 0.0000 103.3870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.1870 0.0000 103.3870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.1870 0.0000 103.3870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.4590 0.0000 74.6590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.4590 0.0000 74.6590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.4590 0.0000 74.6590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.4590 0.0000 74.6590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.4590 0.0000 74.6590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.8270 0.0000 76.0270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.8270 0.0000 76.0270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.8270 0.0000 76.0270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.8270 0.0000 76.0270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.8270 0.0000 76.0270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.1440 0.0000 75.3440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.1440 0.0000 75.3440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.1440 0.0000 75.3440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.1440 0.0000 75.3440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.1440 0.0000 75.3440 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[28]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.5040 0.0000 102.7040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.5040 0.0000 102.7040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.5040 0.0000 102.7040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.5040 0.0000 102.7040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.5040 0.0000 102.7040 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[22]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.6160 0.0000 80.8160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.6160 0.0000 80.8160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.6160 0.0000 80.8160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.6160 0.0000 80.8160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.6160 0.0000 80.8160 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[14]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.6670 0.0000 82.8670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.6670 0.0000 82.8670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.6670 0.0000 82.8670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.6670 0.0000 82.8670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.6670 0.0000 82.8670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.9840 0.0000 82.1840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.9840 0.0000 82.1840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.9840 0.0000 82.1840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.9840 0.0000 82.1840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.9840 0.0000 82.1840 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[6]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 123.7070 0.0000 123.9070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.7070 0.0000 123.9070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.7070 0.0000 123.9070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.7070 0.0000 123.9070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.7070 0.0000 123.9070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 123.0240 0.0000 123.2240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.0240 0.0000 123.2240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.0240 0.0000 123.2240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.0240 0.0000 123.2240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.0240 0.0000 123.2240 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[42]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 118.2350 0.0000 118.4350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.2350 0.0000 118.4350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.2350 0.0000 118.4350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 118.2350 0.0000 118.4350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.2350 0.0000 118.4350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 117.5520 0.0000 117.7520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.5520 0.0000 117.7520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.5520 0.0000 117.7520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 117.5520 0.0000 117.7520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.5520 0.0000 117.7520 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[8]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.9710 0.0000 121.1710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.9710 0.0000 121.1710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.9710 0.0000 121.1710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.9710 0.0000 121.1710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.9710 0.0000 121.1710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.8240 0.0000 89.0240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.8240 0.0000 89.0240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.8240 0.0000 89.0240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.8240 0.0000 89.0240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.8240 0.0000 89.0240 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[10]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.2430 0.0000 92.4430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.2430 0.0000 92.4430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.2430 0.0000 92.4430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.2430 0.0000 92.4430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.2430 0.0000 92.4430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.5600 0.0000 91.7600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.5600 0.0000 91.7600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.5600 0.0000 91.7600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.5600 0.0000 91.7600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.5600 0.0000 91.7600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[25]
  OBS
    LAYER M2 ;
      RECT 0.0000 218.2300 147.6070 219.8200 ;
      RECT 0.0000 212.6000 147.6070 219.8200 ;
      RECT 0.0000 212.6000 148.4910 218.2300 ;
      RECT 0.0000 211.0000 147.5920 212.6000 ;
      RECT 0.0000 209.4100 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 203.7800 148.4910 209.4100 ;
      RECT 0.0000 202.1900 147.5940 203.7800 ;
      RECT 0.0000 200.5900 147.5910 202.1900 ;
      RECT 0.0000 50.7360 148.4910 200.5900 ;
      RECT 0.0000 49.1360 147.5910 50.7360 ;
      RECT 0.0000 18.1900 148.4910 49.1360 ;
      RECT 0.0000 16.1280 147.5910 18.1900 ;
      RECT 0.0000 10.7180 148.4910 16.1280 ;
      RECT 0.0000 9.1180 147.5910 10.7180 ;
      RECT 0.0000 0.9000 148.4910 9.1180 ;
      RECT 0.0000 0.0000 64.1830 0.9000 ;
      RECT 128.7000 0.0000 148.4910 9.1180 ;
      RECT 128.7000 0.0000 148.4910 0.9000 ;
      RECT 0.0000 247.8670 148.4910 264.7580 ;
      RECT 0.0000 228.6500 147.5970 264.7580 ;
      RECT 0.0000 0.0000 64.1830 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 242.8910 147.5970 247.8670 ;
      RECT 0.0000 228.6500 148.4910 242.8910 ;
      RECT 0.0000 227.0500 147.5910 228.6500 ;
      RECT 147.5970 245.1150 148.4910 246.2670 ;
      RECT 0.0000 221.4200 148.4910 227.0500 ;
      RECT 0.0000 212.6000 147.5940 227.0500 ;
      RECT 0.0000 202.1900 147.5920 227.0500 ;
      RECT 0.0000 219.8200 147.5940 221.4200 ;
    LAYER M1 ;
      RECT 147.7070 219.7300 148.4910 219.9200 ;
      RECT 147.6940 202.0900 148.4910 202.2800 ;
      RECT 147.6940 210.9100 148.4910 211.1000 ;
      RECT 147.6970 245.0150 148.4910 246.3670 ;
      RECT 0.0000 221.3200 148.4910 227.1500 ;
      RECT 0.0000 212.5000 147.6940 227.1500 ;
      RECT 0.0000 202.0900 147.6920 227.1500 ;
      RECT 0.0000 219.9200 147.6940 221.3200 ;
      RECT 0.0000 218.3300 147.7070 219.9200 ;
      RECT 0.0000 212.5000 147.7070 219.9200 ;
      RECT 0.0000 212.5000 148.4910 218.3300 ;
      RECT 0.0000 211.1000 147.6920 212.5000 ;
      RECT 0.0000 209.5100 147.6940 211.1000 ;
      RECT 0.0000 202.0900 147.6940 211.1000 ;
      RECT 0.0000 202.0900 147.6940 211.1000 ;
      RECT 0.0000 203.6800 148.4910 209.5100 ;
      RECT 0.0000 202.0900 147.6940 203.6800 ;
      RECT 0.0000 200.6900 147.6910 202.0900 ;
      RECT 0.0000 50.6360 148.4910 200.6900 ;
      RECT 0.0000 49.2360 147.6910 50.6360 ;
      RECT 0.0000 18.0900 148.4910 49.2360 ;
      RECT 0.0000 16.2280 147.6910 18.0900 ;
      RECT 0.0000 10.6180 148.4910 16.2280 ;
      RECT 0.0000 9.2180 147.6910 10.6180 ;
      RECT 0.0000 0.8000 148.4910 9.2180 ;
      RECT 0.0000 0.0000 64.2830 0.8000 ;
      RECT 128.6000 0.0000 148.4910 9.2180 ;
      RECT 128.6000 0.0000 148.4910 0.8000 ;
      RECT 0.0000 247.7670 148.4910 264.7580 ;
      RECT 0.0000 228.5500 147.6970 264.7580 ;
      RECT 0.0000 0.0000 64.2830 264.7580 ;
      RECT 0.0000 0.8000 147.6910 264.7580 ;
      RECT 0.0000 0.8000 147.6910 264.7580 ;
      RECT 0.0000 0.8000 147.6910 264.7580 ;
      RECT 0.0000 0.8000 147.6910 264.7580 ;
      RECT 0.0000 0.8000 147.6910 264.7580 ;
      RECT 0.0000 242.9910 147.6970 247.7670 ;
      RECT 0.0000 228.5500 148.4910 242.9910 ;
      RECT 0.0000 227.1500 147.6910 228.5500 ;
    LAYER PO ;
      RECT 0.0000 0.0000 148.4910 264.7580 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 148.4910 264.7580 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 148.4910 264.7580 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 148.4910 264.7580 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 148.4910 264.7580 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 148.4910 264.7580 ;
    LAYER M5 ;
      RECT 148.1500 263.7570 148.4910 264.7580 ;
      RECT 147.5970 245.1150 148.4910 246.2670 ;
      RECT 0.0000 0.0000 64.1830 0.9000 ;
      RECT 128.7000 0.0000 148.4910 0.9000 ;
      RECT 0.0000 263.7570 144.6500 263.7580 ;
      RECT 0.0000 0.9000 65.5510 263.7580 ;
      RECT 0.0000 0.9010 144.6500 263.7580 ;
      RECT 0.0000 247.8670 148.4910 263.7570 ;
      RECT 0.0000 228.6500 147.5970 263.7570 ;
      RECT 0.0000 0.9010 147.5910 263.7570 ;
      RECT 0.0000 0.9010 147.5910 263.7570 ;
      RECT 0.0000 0.9010 147.5910 263.7570 ;
      RECT 0.0000 0.9010 147.5910 263.7570 ;
      RECT 0.0000 0.9010 147.5910 263.7570 ;
      RECT 0.0000 242.8910 147.5970 247.8670 ;
      RECT 0.0000 228.6500 148.4910 242.8910 ;
      RECT 0.0000 227.0500 147.5910 228.6500 ;
      RECT 0.0000 221.4200 148.4910 227.0500 ;
      RECT 0.0000 212.6000 147.5940 227.0500 ;
      RECT 0.0000 202.1900 147.5920 227.0500 ;
      RECT 0.0000 219.8200 147.5940 221.4200 ;
      RECT 0.0000 218.2300 147.6070 219.8200 ;
      RECT 0.0000 212.6000 147.6070 219.8200 ;
      RECT 0.0000 212.6000 148.4910 218.2300 ;
      RECT 0.0000 211.0000 147.5920 212.6000 ;
      RECT 0.0000 209.4100 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 203.7800 148.4910 209.4100 ;
      RECT 0.0000 202.1900 147.5940 203.7800 ;
      RECT 0.0000 200.5900 147.5910 202.1900 ;
      RECT 0.0000 50.7360 148.4910 200.5900 ;
      RECT 0.0000 49.1360 147.5910 50.7360 ;
      RECT 0.0000 18.1900 148.4910 49.1360 ;
      RECT 0.0000 16.1280 147.5910 18.1900 ;
      RECT 0.0000 10.7180 148.4910 16.1280 ;
      RECT 0.0000 9.1180 147.5910 10.7180 ;
      RECT 0.0000 0.9010 148.4910 9.1180 ;
      RECT 0.0000 0.9000 65.5510 0.9010 ;
      RECT 67.1510 0.9000 148.4910 9.1180 ;
      RECT 67.1510 0.9000 148.4910 0.9010 ;
      RECT 128.7000 0.0000 148.4910 9.1180 ;
    LAYER M4 ;
      RECT 147.5970 245.1150 148.4910 246.2670 ;
      RECT 128.7000 0.0000 148.4910 0.9000 ;
      RECT 0.0000 0.0000 64.1830 0.9000 ;
      RECT 0.0000 221.4200 148.4910 227.0500 ;
      RECT 0.0000 212.6000 147.5940 227.0500 ;
      RECT 0.0000 202.1900 147.5920 227.0500 ;
      RECT 0.0000 219.8200 147.5940 221.4200 ;
      RECT 0.0000 218.2300 147.6070 219.8200 ;
      RECT 0.0000 212.6000 147.6070 219.8200 ;
      RECT 0.0000 212.6000 148.4910 218.2300 ;
      RECT 0.0000 211.0000 147.5920 212.6000 ;
      RECT 0.0000 209.4100 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 203.7800 148.4910 209.4100 ;
      RECT 0.0000 202.1900 147.5940 203.7800 ;
      RECT 0.0000 200.5900 147.5910 202.1900 ;
      RECT 0.0000 50.7360 148.4910 200.5900 ;
      RECT 0.0000 49.1360 147.5910 50.7360 ;
      RECT 0.0000 18.1900 148.4910 49.1360 ;
      RECT 0.0000 16.1280 147.5910 18.1900 ;
      RECT 0.0000 10.7180 148.4910 16.1280 ;
      RECT 0.0000 9.1180 147.5910 10.7180 ;
      RECT 0.0000 0.9010 148.4910 9.1180 ;
      RECT 0.0000 0.9000 65.5510 0.9010 ;
      RECT 67.1510 0.9000 148.4910 9.1180 ;
      RECT 67.1510 0.9000 148.4910 0.9010 ;
      RECT 0.0000 247.8670 148.4910 264.7580 ;
      RECT 0.0000 228.6500 147.5970 264.7580 ;
      RECT 0.0000 0.0000 64.1830 264.7580 ;
      RECT 0.0000 0.9000 65.5510 264.7580 ;
      RECT 0.0000 0.9010 147.5910 264.7580 ;
      RECT 0.0000 0.9010 147.5910 264.7580 ;
      RECT 0.0000 0.9010 147.5910 264.7580 ;
      RECT 0.0000 0.9010 147.5910 264.7580 ;
      RECT 0.0000 0.9010 147.5910 264.7580 ;
      RECT 0.0000 242.8910 147.5970 247.8670 ;
      RECT 0.0000 228.6500 148.4910 242.8910 ;
      RECT 0.0000 227.0500 147.5910 228.6500 ;
    LAYER M3 ;
      RECT 147.5970 245.1150 148.4910 246.2670 ;
      RECT 0.0000 221.4200 148.4910 227.0500 ;
      RECT 0.0000 212.6000 147.5940 227.0500 ;
      RECT 0.0000 202.1900 147.5920 227.0500 ;
      RECT 0.0000 219.8200 147.5940 221.4200 ;
      RECT 0.0000 218.2300 147.6070 219.8200 ;
      RECT 0.0000 212.6000 147.6070 219.8200 ;
      RECT 0.0000 212.6000 148.4910 218.2300 ;
      RECT 0.0000 211.0000 147.5920 212.6000 ;
      RECT 0.0000 209.4100 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 202.1900 147.5940 211.0000 ;
      RECT 0.0000 203.7800 148.4910 209.4100 ;
      RECT 0.0000 202.1900 147.5940 203.7800 ;
      RECT 0.0000 200.5900 147.5910 202.1900 ;
      RECT 0.0000 50.7360 148.4910 200.5900 ;
      RECT 0.0000 49.1360 147.5910 50.7360 ;
      RECT 0.0000 18.1900 148.4910 49.1360 ;
      RECT 0.0000 16.1280 147.5910 18.1900 ;
      RECT 0.0000 10.7180 148.4910 16.1280 ;
      RECT 0.0000 9.1180 147.5910 10.7180 ;
      RECT 0.0000 0.9000 148.4910 9.1180 ;
      RECT 0.0000 0.0000 64.1830 0.9000 ;
      RECT 128.7000 0.0000 148.4910 9.1180 ;
      RECT 128.7000 0.0000 148.4910 0.9000 ;
      RECT 0.0000 247.8670 148.4910 264.7580 ;
      RECT 0.0000 228.6500 147.5970 264.7580 ;
      RECT 0.0000 0.0000 64.1830 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 0.9000 147.5910 264.7580 ;
      RECT 0.0000 242.8910 147.5970 247.8670 ;
      RECT 0.0000 228.6500 148.4910 242.8910 ;
      RECT 0.0000 227.0500 147.5910 228.6500 ;
  END
END SRAMLP1RW256x46

MACRO SRAMLP1RW256x48
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 155.143 BY 268.197 ;
  SYMMETRY X Y R90 ;

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.3500 0.0000 76.5500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.3500 0.0000 76.5500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.3500 0.0000 76.5500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.3500 0.0000 76.5500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.3500 0.0000 76.5500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[7]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.5470 0.0000 110.7470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.5470 0.0000 110.7470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.5470 0.0000 110.7470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.5470 0.0000 110.7470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.5470 0.0000 110.7470 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[30]

  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.2370 0.0000 98.4370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.2370 0.0000 98.4370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.2370 0.0000 98.4370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.2370 0.0000 98.4370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.2370 0.0000 98.4370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[46]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.9830 0.0000 75.1830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.9830 0.0000 75.1830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.9830 0.0000 75.1830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.9830 0.0000 75.1830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.9830 0.0000 75.1830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[6]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.9240 0.0000 86.1240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.9240 0.0000 86.1240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.9240 0.0000 86.1240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.9240 0.0000 86.1240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.9240 0.0000 86.1240 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M2 ;
  END O[13]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.6120 0.0000 73.8120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.6120 0.0000 73.8120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.6120 0.0000 73.8120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.6120 0.0000 73.8120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.6120 0.0000 73.8120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[4]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.7260 0.0000 77.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.7260 0.0000 77.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.7260 0.0000 77.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.7260 0.0000 77.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.7260 0.0000 77.9260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[8]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.2460 0.0000 72.4460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.2460 0.0000 72.4460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.2460 0.0000 72.4460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.2460 0.0000 72.4460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.2460 0.0000 72.4460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1412 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1412 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1412 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1412 LAYER M2 ;
  END O[1]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.8770 0.0000 71.0770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.8770 0.0000 71.0770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.8770 0.0000 71.0770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.8770 0.0000 71.0770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.8770 0.0000 71.0770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[0]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.2940 0.0000 87.4940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.2940 0.0000 87.4940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.2940 0.0000 87.4940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.2940 0.0000 87.4940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.2940 0.0000 87.4940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[14]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.6610 0.0000 88.8610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.6610 0.0000 88.8610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.6610 0.0000 88.8610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.6610 0.0000 88.8610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.6610 0.0000 88.8610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[15]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.0920 0.0000 79.2920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.0920 0.0000 79.2920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.0920 0.0000 79.2920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.0920 0.0000 79.2920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.0920 0.0000 79.2920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[9]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.5560 0.0000 84.7560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.5560 0.0000 84.7560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.5560 0.0000 84.7560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.5560 0.0000 84.7560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.5560 0.0000 84.7560 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[12]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.8230 0.0000 82.0230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.8230 0.0000 82.0230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.8230 0.0000 82.0230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.8230 0.0000 82.0230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.8230 0.0000 82.0230 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[11]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 114.6460 0.0000 114.8460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.6460 0.0000 114.8460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.6460 0.0000 114.8460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.6460 0.0000 114.8460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.6460 0.0000 114.8460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[32]

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 113.2810 0.0000 113.4810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.2810 0.0000 113.4810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.2810 0.0000 113.4810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 113.2810 0.0000 113.4810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.2810 0.0000 113.4810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[45]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.9110 0.0000 112.1110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.9110 0.0000 112.1110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.9110 0.0000 112.1110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.9110 0.0000 112.1110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.9110 0.0000 112.1110 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[31]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.1420 0.0000 68.3420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.1420 0.0000 68.3420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.1420 0.0000 68.3420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.1420 0.0000 68.3420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.1420 0.0000 68.3420 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[42]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 130.4110 0.0000 130.6110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.4110 0.0000 130.6110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.4110 0.0000 130.6110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 130.4110 0.0000 130.6110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 130.4110 0.0000 130.6110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9490 256.0990 155.1430 256.2990 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9490 256.0990 155.1430 256.2990 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9490 256.0990 155.1430 256.2990 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9490 256.0990 155.1430 256.2990 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9490 256.0990 155.1430 256.2990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.7780 0.0000 131.9780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.7780 0.0000 131.9780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.7780 0.0000 131.9780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.7780 0.0000 131.9780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.7780 0.0000 131.9780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9490 257.2600 155.1430 257.4600 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9490 257.2600 155.1430 257.4600 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9490 257.2600 155.1430 257.4600 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9490 257.2600 155.1430 257.4600 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9490 257.2600 155.1430 257.4600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.3950 0.0000 91.5950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.3950 0.0000 91.5950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.3950 0.0000 91.5950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.3950 0.0000 91.5950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.3950 0.0000 91.5950 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[17]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.0300 0.0000 90.2300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.0300 0.0000 90.2300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.0300 0.0000 90.2300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.0300 0.0000 90.2300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.0300 0.0000 90.2300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[16]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.5020 0.0000 95.7020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.5020 0.0000 95.7020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.5020 0.0000 95.7020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.5020 0.0000 95.7020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.5020 0.0000 95.7020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[20]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.1300 0.0000 94.3300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.1300 0.0000 94.3300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.1300 0.0000 94.3300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.1300 0.0000 94.3300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.1300 0.0000 94.3300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[19]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.7730 0.0000 92.9730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.7730 0.0000 92.9730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.7730 0.0000 92.9730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.7730 0.0000 92.9730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.7730 0.0000 92.9730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[18]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.6050 0.0000 99.8050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.6050 0.0000 99.8050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.6050 0.0000 99.8050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.6050 0.0000 99.8050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.6050 0.0000 99.8050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[22]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.4610 0.0000 80.6610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.4610 0.0000 80.6610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.4610 0.0000 80.6610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.4610 0.0000 80.6610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.4610 0.0000 80.6610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[10]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.8700 0.0000 97.0700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.8700 0.0000 97.0700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.8700 0.0000 97.0700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.8700 0.0000 97.0700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.8700 0.0000 97.0700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[21]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.7090 0.0000 103.9090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.7090 0.0000 103.9090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.7090 0.0000 103.9090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.7090 0.0000 103.9090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.7090 0.0000 103.9090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[25]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.3410 0.0000 102.5410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.3410 0.0000 102.5410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.3410 0.0000 102.5410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.3410 0.0000 102.5410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.3410 0.0000 102.5410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[24]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.9730 0.0000 101.1730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.9730 0.0000 101.1730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.9730 0.0000 101.1730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.9730 0.0000 101.1730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.9730 0.0000 101.1730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[23]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.4480 0.0000 106.6480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.4480 0.0000 106.6480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.4480 0.0000 106.6480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.4480 0.0000 106.6480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.4480 0.0000 106.6480 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[27]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.0740 0.0000 105.2740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.0740 0.0000 105.2740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.0740 0.0000 105.2740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.0740 0.0000 105.2740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.0740 0.0000 105.2740 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[26]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.8130 0.0000 108.0130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.8130 0.0000 108.0130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.8140 0.0000 108.0140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.8140 0.0000 108.0140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.8140 0.0000 108.0140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[28]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.4750 0.0000 67.6750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.4750 0.0000 67.6750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.4750 0.0000 67.6750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.4750 0.0000 67.6750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.4750 0.0000 67.6750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[42]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8430 0.0000 69.0430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8430 0.0000 69.0430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8430 0.0000 69.0430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8430 0.0000 69.0430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8430 0.0000 69.0430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.5730 0.0000 97.7730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.5730 0.0000 97.7730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.5730 0.0000 97.7730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.5730 0.0000 97.7730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.5730 0.0000 97.7730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[46]

  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.5230 0.0000 82.7230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.5230 0.0000 82.7230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.5230 0.0000 82.7230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.5230 0.0000 82.7230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.5230 0.0000 82.7230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[47]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.7290 0.0000 116.9290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.7290 0.0000 116.9290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.7290 0.0000 116.9290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.7290 0.0000 116.9290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.7290 0.0000 116.9290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 118.0990 0.0000 118.2990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.0990 0.0000 118.2990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.0990 0.0000 118.2990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 118.0990 0.0000 118.2990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.0990 0.0000 118.2990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 119.4640 0.0000 119.6640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.4640 0.0000 119.6640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.4640 0.0000 119.6640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.4640 0.0000 119.6640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.4640 0.0000 119.6640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.8330 0.0000 121.0330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.8330 0.0000 121.0330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.8330 0.0000 121.0330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.8330 0.0000 121.0330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.8330 0.0000 121.0330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 122.2030 0.0000 122.4030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.2030 0.0000 122.4030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.2030 0.0000 122.4030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 122.2030 0.0000 122.4030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.2030 0.0000 122.4030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[37]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 123.5680 0.0000 123.7680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.5680 0.0000 123.7680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.5680 0.0000 123.7680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.5680 0.0000 123.7680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.5680 0.0000 123.7680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 124.9350 0.0000 125.1350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.9350 0.0000 125.1350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.9350 0.0000 125.1350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 124.9350 0.0000 125.1350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.9350 0.0000 125.1350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[39]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 126.3060 0.0000 126.5060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.3060 0.0000 126.5060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.3060 0.0000 126.5060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 126.3060 0.0000 126.5060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 126.3060 0.0000 126.5060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[40]

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 50.9100 155.1430 51.1100 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 50.9100 155.1430 51.1100 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 50.9100 155.1430 51.1100 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 50.9100 155.1430 51.1100 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 50.9100 155.1430 51.1100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 127.6730 0.0000 127.8730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.6730 0.0000 127.8730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.6730 0.0000 127.8730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 127.6730 0.0000 127.8730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 127.6730 0.0000 127.8730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[41]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 133.1390 0.0000 133.3390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.1390 0.0000 133.3390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.1390 0.0000 133.3390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 133.1390 0.0000 133.3390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 133.1390 0.0000 133.3390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 129.0390 0.0000 129.2390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.0390 0.0000 129.2390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.0390 0.0000 129.2390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.0390 0.0000 129.2390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 129.0390 0.0000 129.2390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 16.8340 155.1430 17.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 16.8340 155.1430 17.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 16.8340 155.1430 17.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 16.8340 155.1430 17.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 16.8340 155.1430 17.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.6830 0.0000 75.8830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.6830 0.0000 75.8830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.6830 0.0000 75.8830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.6830 0.0000 75.8830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.6830 0.0000 75.8830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 115.3590 0.0000 115.5590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.3590 0.0000 115.5590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.3590 0.0000 115.5590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.3590 0.0000 115.5590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.3590 0.0000 115.5590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.8840 0.0000 110.0840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.8840 0.0000 110.0840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.8840 0.0000 110.0840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.8840 0.0000 110.0840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.8840 0.0000 110.0840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.2130 0.0000 70.4130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.2130 0.0000 70.4130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.2130 0.0000 70.4130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.2130 0.0000 70.4130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.2130 0.0000 70.4130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.3140 0.0000 74.5140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.3140 0.0000 74.5140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.3140 0.0000 74.5140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.3140 0.0000 74.5140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.3140 0.0000 74.5140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.2600 0.0000 85.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.2600 0.0000 85.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.2600 0.0000 85.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.2600 0.0000 85.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.2600 0.0000 85.4600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.9460 0.0000 73.1460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.9460 0.0000 73.1460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.9460 0.0000 73.1460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.9460 0.0000 73.1460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.9460 0.0000 73.1460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.4280 0.0000 78.6280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.4280 0.0000 78.6280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.4280 0.0000 78.6280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.4280 0.0000 78.6280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.4280 0.0000 78.6280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.6220 0.0000 86.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.6220 0.0000 86.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.6220 0.0000 86.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.6220 0.0000 86.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.6220 0.0000 86.8220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.0500 0.0000 77.2500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.0500 0.0000 77.2500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.0500 0.0000 77.2500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.0500 0.0000 77.2500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.0500 0.0000 77.2500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.5780 0.0000 71.7780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.5780 0.0000 71.7780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.5780 0.0000 71.7780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.5780 0.0000 71.7780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.5780 0.0000 71.7780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.1560 0.0000 81.3560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.1560 0.0000 81.3560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.1560 0.0000 81.3560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.1560 0.0000 81.3560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.1560 0.0000 81.3560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9940 0.0000 88.1940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9940 0.0000 88.1940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9940 0.0000 88.1940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9940 0.0000 88.1940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9940 0.0000 88.1940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 2.8240 267.8970 3.1240 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.7240 267.8970 4.0240 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.9070 267.8970 128.2070 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.8070 267.8970 129.1070 268.1970 ;
    END
  END VDDL

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 113.9960 0.0000 114.1960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.9960 0.0000 114.1960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.9960 0.0000 114.1960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 113.9960 0.0000 114.1960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.9960 0.0000 114.1960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.8910 0.0000 84.0910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.8910 0.0000 84.0910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.8910 0.0000 84.0910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.8910 0.0000 84.0910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.8910 0.0000 84.0910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 112.6260 0.0000 112.8260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.6260 0.0000 112.8260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.6260 0.0000 112.8260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 112.6260 0.0000 112.8260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.6260 0.0000 112.8260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.2520 0.0000 111.4520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.2520 0.0000 111.4520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.2520 0.0000 111.4520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.2520 0.0000 111.4520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.2520 0.0000 111.4520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.3080 0.0000 100.5080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.3080 0.0000 100.5080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.3080 0.0000 100.5080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.3080 0.0000 100.5080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.3080 0.0000 100.5080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 219.7960 155.1430 219.9960 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 219.7960 155.1430 219.9960 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 219.7960 155.1430 219.9960 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 219.7960 155.1430 219.9960 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 219.7960 155.1430 219.9960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.23404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23404 LAYER M3 ;
    ANTENNAMAXAREACAR 22.9276 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 27.06817 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 31.20846 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[2]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 229.0720 155.1430 229.2720 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 229.0720 155.1430 229.2720 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 229.0720 155.1430 229.2720 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 229.0720 155.1430 229.2720 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 229.0720 155.1430 229.2720 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2365 LAYER M3 ;
    ANTENNAMAXAREACAR 22.98776 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 27.12832 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 31.26861 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[0]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9490 260.6300 155.1430 260.8300 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9490 260.6300 155.1430 260.8300 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9490 260.6300 155.1430 260.8300 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9490 260.6300 155.1430 260.8300 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9490 260.6300 155.1430 260.8300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 2.3406 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 5.563501 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 5.563501 LAYER M1 ;
    ANTENNAGATEAREA 2.3406 LAYER M2 ;
    ANTENNAGATEAREA 2.3406 LAYER M3 ;
    ANTENNAGATEAREA 2.3406 LAYER M4 ;
    ANTENNAGATEAREA 2.3406 LAYER M5 ;
    ANTENNAGATEAREA 2.3406 LAYER M6 ;
    ANTENNAGATEAREA 2.3406 LAYER M7 ;
    ANTENNAGATEAREA 2.3406 LAYER M8 ;
    ANTENNAGATEAREA 2.3406 LAYER M9 ;
    ANTENNAGATEAREA 2.3406 LAYER MRDL ;
  END LS

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 202.9860 155.1430 203.1860 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 202.9860 155.1430 203.1860 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 202.9860 155.1430 203.1860 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 202.9860 155.1430 203.1860 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 202.9860 155.1430 203.1860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.183 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 7.620792 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 7.620792 LAYER M1 ;
    ANTENNAGATEAREA 68.6994 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 6441.221 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6441.221 LAYER M2 ;
    ANTENNAMAXAREACAR 213.9628 LAYER M2 ;
    ANTENNAGATEAREA 81.6288 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 927.1143 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 927.1143 LAYER M3 ;
    ANTENNAMAXAREACAR 742.8267 LAYER M3 ;
    ANTENNAGATEAREA 81.6288 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 5730.405 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5730.405 LAYER M4 ;
    ANTENNAMAXAREACAR 813.0275 LAYER M4 ;
    ANTENNAGATEAREA 81.6288 LAYER M5 ;
    ANTENNAGATEAREA 81.6288 LAYER M6 ;
    ANTENNAGATEAREA 81.6288 LAYER M7 ;
    ANTENNAGATEAREA 81.6288 LAYER M8 ;
    ANTENNAGATEAREA 81.6288 LAYER M9 ;
    ANTENNAGATEAREA 81.6288 LAYER MRDL ;
  END A[5]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.1000 0.0000 92.3000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.1000 0.0000 92.3000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.1000 0.0000 92.3000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.1000 0.0000 92.3000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.1000 0.0000 92.3000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.3650 0.0000 89.5650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.3650 0.0000 89.5650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.3650 0.0000 89.5650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.3650 0.0000 89.5650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.3650 0.0000 89.5650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.7330 0.0000 90.9330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.7330 0.0000 90.9330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.7330 0.0000 90.9330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.7330 0.0000 90.9330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.7330 0.0000 90.9330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.2050 0.0000 96.4050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.2050 0.0000 96.4050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.2050 0.0000 96.4050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.2050 0.0000 96.4050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.2050 0.0000 96.4050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.8350 0.0000 95.0350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.8350 0.0000 95.0350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.8350 0.0000 95.0350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.8350 0.0000 95.0350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.8350 0.0000 95.0350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.4670 0.0000 93.6670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.4670 0.0000 93.6670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.4670 0.0000 93.6670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.4670 0.0000 93.6670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.4670 0.0000 93.6670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.9380 0.0000 99.1380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.9380 0.0000 99.1380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.9380 0.0000 99.1380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.9380 0.0000 99.1380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.9380 0.0000 99.1380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.7860 0.0000 79.9860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.7860 0.0000 79.9860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.7860 0.0000 79.9860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.7860 0.0000 79.9860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.7860 0.0000 79.9860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.4110 0.0000 104.6110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.4110 0.0000 104.6110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.4110 0.0000 104.6110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.4110 0.0000 104.6110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.4110 0.0000 104.6110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.0430 0.0000 103.2430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.0430 0.0000 103.2430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.0430 0.0000 103.2430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.0430 0.0000 103.2430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.0430 0.0000 103.2430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.6750 0.0000 101.8750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.6750 0.0000 101.8750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.6750 0.0000 101.8750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.6750 0.0000 101.8750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.6750 0.0000 101.8750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.1470 0.0000 107.3470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.1470 0.0000 107.3470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.1470 0.0000 107.3470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.1470 0.0000 107.3470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.1470 0.0000 107.3470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.7790 0.0000 105.9790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.7790 0.0000 105.9790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.7790 0.0000 105.9790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.7790 0.0000 105.9790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.7790 0.0000 105.9790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.5150 0.0000 108.7150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.5150 0.0000 108.7150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.5150 0.0000 108.7150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.5150 0.0000 108.7150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.5150 0.0000 108.7150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 1.0240 267.8970 1.3230 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9250 267.8970 2.2260 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.7080 267.8970 130.0080 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.6070 267.8970 130.9060 268.1970 ;
    END
  END VDD

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 220.5250 155.1430 220.7250 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 220.5250 155.1430 220.7250 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 220.5250 155.1430 220.7250 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 220.5250 155.1430 220.7250 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 220.5250 155.1430 220.7250 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.23866 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23866 LAYER M3 ;
    ANTENNAMAXAREACAR 24.67288 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 28.81333 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 32.9535 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[1]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 202.3650 155.1430 202.5650 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 202.3650 155.1430 202.5650 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 202.3650 155.1430 202.5650 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 202.3650 155.1430 202.5650 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 202.3650 155.1430 202.5650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.784278 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.784278 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAMAXAREACAR 25.56902 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 29.70941 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 33.84953 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 37.98937 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[6]

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 3.2740 267.8970 3.5730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.1750 267.8970 4.4760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4740 267.8970 1.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3750 267.8970 2.6750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.5740 267.8970 0.8740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8750 267.8970 7.1750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7740 267.8970 8.0730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6750 267.8970 8.9760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0740 267.8970 5.3740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9740 267.8970 6.2740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0740 267.8970 14.3740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1740 267.8970 13.4740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2740 267.8970 12.5740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4740 267.8970 10.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3750 267.8970 11.6750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5740 267.8970 9.8740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6740 267.8970 17.9740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7740 267.8970 17.0740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8740 267.8970 16.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5750 267.8970 18.8750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9750 267.8970 15.2750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0730 267.8970 23.3730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2730 267.8970 21.5730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3740 267.8970 20.6740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4740 267.8970 19.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1740 267.8970 22.4740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7750 267.8970 26.0740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9750 267.8970 24.2750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8750 267.8970 25.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6740 267.8970 26.9750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5740 267.8970 27.8750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4740 267.8970 28.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2750 267.8970 30.5750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9740 267.8970 33.2740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0750 267.8970 32.3760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3740 267.8970 29.6740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1740 267.8970 31.4730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4740 267.8970 37.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6740 267.8970 35.9730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5750 267.8970 36.8760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8740 267.8970 34.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7750 267.8970 35.0750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2750 267.8970 39.5750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1740 267.8970 40.4730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0750 267.8970 41.3760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3740 267.8970 38.6740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8740 267.8970 43.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9740 267.8970 42.2740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4740 267.8970 46.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5740 267.8970 45.8740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6740 267.8970 44.9740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3750 267.8970 47.6750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7750 267.8970 44.0750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8740 267.8970 52.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0740 267.8970 50.3740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1740 267.8970 49.4740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2740 267.8970 48.5740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9750 267.8970 51.2750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3750 267.8970 56.6750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2750 267.8970 57.5740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4730 267.8970 55.7730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6730 267.8970 53.9730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7740 267.8970 53.0740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5740 267.8970 54.8740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0740 267.8970 59.3750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9740 267.8970 60.2750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7740 267.8970 62.0740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8740 267.8970 61.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1750 267.8970 58.4740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2740 267.8970 66.5740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6750 267.8970 62.9750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3740 267.8970 65.6740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4750 267.8970 64.7760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5740 267.8970 63.8730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6750 267.8970 71.9750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8740 267.8970 70.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0740 267.8970 68.3730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9750 267.8970 69.2760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1750 267.8970 67.4750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7740 267.8970 71.0740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5740 267.8970 72.8730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4750 267.8970 73.7760 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2740 267.8970 75.5740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1750 267.8970 76.4750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3740 267.8970 74.6740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5740 267.8970 81.8740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6740 267.8970 80.9740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8740 267.8970 79.1740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9740 267.8970 78.2740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.0740 267.8970 77.3740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7750 267.8970 80.0750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0730 267.8970 86.3730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1740 267.8970 85.4740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2740 267.8970 84.5740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4740 267.8970 82.7740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3750 267.8970 83.6750 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.7600 267.8970 89.0600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.6600 267.8970 89.9590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.8730 267.8970 88.1730 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.9740 267.8970 87.2740 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.5600 267.8970 90.8590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.0600 267.8970 95.3600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.4590 267.8970 91.7600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.3590 267.8970 92.6600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.1590 267.8970 94.4590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.2590 267.8970 93.5590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.9590 267.8970 96.2580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.4590 267.8970 100.7580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.6590 267.8970 98.9590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.5600 267.8970 99.8600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.7590 267.8970 98.0590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.8600 267.8970 97.1610 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.0600 267.8970 104.3600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.9590 267.8970 105.2580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.2590 267.8970 102.5590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.3600 267.8970 101.6610 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.1590 267.8970 103.4590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.8600 267.8970 106.1610 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.3590 267.8970 110.6590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.4590 267.8970 109.7590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.6590 267.8970 107.9590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.5600 267.8970 108.8600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.7590 267.8970 107.0590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.8590 267.8970 115.1590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.9590 267.8970 114.2590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.0590 267.8970 113.3590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.2590 267.8970 111.5590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.1600 267.8970 112.4600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.4580 267.8970 118.7580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.5590 267.8970 117.8590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.6590 267.8970 116.9590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.3590 267.8970 119.6590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.7600 267.8970 116.0600 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.1580 267.8970 121.4580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.0580 267.8970 122.3570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.8570 267.8970 124.1580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.7570 267.8970 125.0580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.2580 267.8970 120.5580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.9580 267.8970 123.2570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.4580 267.8970 127.7580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.2580 267.8970 129.5590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.5570 267.8970 126.8570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.6570 267.8970 125.9570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.3570 267.8970 128.6560 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.8570 267.8970 133.1560 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.7580 267.8970 134.0590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.0570 267.8970 131.3570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.9580 267.8970 132.2580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.1570 267.8970 130.4570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.4580 267.8970 136.7580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.3570 267.8970 137.6560 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.2580 267.8970 138.5590 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.6570 267.8970 134.9570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.5570 267.8970 135.8570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.1570 267.8970 139.4570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.6570 267.8970 143.9570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.7570 267.8970 143.0570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.8570 267.8970 142.1570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.0570 267.8970 140.3570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.9580 267.8970 141.2580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.2570 267.8970 147.5570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.3570 267.8970 146.6570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.4570 267.8970 145.7570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.1580 267.8970 148.4580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.7570 267.8970 152.0570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.0570 267.8970 149.3570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.9570 267.8970 150.2570 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.8560 267.8970 151.1560 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.6560 267.8970 152.9560 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.5580 267.8970 153.8580 268.1970 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.5580 267.8970 144.8580 268.1970 ;
    END
  END VSS

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.5120 0.0000 69.7120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.5120 0.0000 69.7120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.5120 0.0000 69.7120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.5120 0.0000 69.7120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.5120 0.0000 69.7120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[44]

  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.1880 0.0000 83.3880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.1880 0.0000 83.3880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.1880 0.0000 83.3880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.1880 0.0000 83.3880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.1880 0.0000 83.3880 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[47]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.0150 0.0000 116.2150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.0150 0.0000 116.2150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.0150 0.0000 116.2150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.0150 0.0000 116.2150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.0150 0.0000 116.2150 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1412 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1412 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1412 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1412 LAYER M2 ;
  END O[33]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 117.3810 0.0000 117.5810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.3810 0.0000 117.5810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.3810 0.0000 117.5810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 117.3810 0.0000 117.5810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.3810 0.0000 117.5810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[34]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 118.7520 0.0000 118.9520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.7520 0.0000 118.9520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.7520 0.0000 118.9520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 118.7520 0.0000 118.9520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.7520 0.0000 118.9520 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[43]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.1190 0.0000 120.3190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.1190 0.0000 120.3190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.1190 0.0000 120.3190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.1190 0.0000 120.3190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.1190 0.0000 120.3190 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[35]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 121.4950 0.0000 121.6950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.4950 0.0000 121.6950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.4950 0.0000 121.6950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 121.4950 0.0000 121.6950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.4950 0.0000 121.6950 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[36]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 122.8610 0.0000 123.0610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.8610 0.0000 123.0610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.8610 0.0000 123.0610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 122.8610 0.0000 123.0610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.8610 0.0000 123.0610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[37]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 124.2300 0.0000 124.4300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.2300 0.0000 124.4300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.2300 0.0000 124.4300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 124.2300 0.0000 124.4300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.2300 0.0000 124.4300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[38]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 125.5920 0.0000 125.7920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.5920 0.0000 125.7920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.5920 0.0000 125.7920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 125.5920 0.0000 125.7920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 125.5920 0.0000 125.7920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[39]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 126.9570 0.0000 127.1570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.9570 0.0000 127.1570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.9570 0.0000 127.1570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 126.9570 0.0000 127.1570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 126.9570 0.0000 127.1570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[40]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 128.3250 0.0000 128.5250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.3250 0.0000 128.5250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.3250 0.0000 128.5250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 128.3250 0.0000 128.5250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 128.3250 0.0000 128.5250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[41]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 129.6930 0.0000 129.8930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.6930 0.0000 129.8930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.6930 0.0000 129.8930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.6930 0.0000 129.8930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 129.6930 0.0000 129.8930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1536 LAYER M2 ;
  END O[2]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.0630 0.0000 131.2630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.0630 0.0000 131.2630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.0630 0.0000 131.2630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.0630 0.0000 131.2630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.0630 0.0000 131.2630 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[3]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.4300 0.0000 132.6300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.4300 0.0000 132.6300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.4300 0.0000 132.6300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.4300 0.0000 132.6300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.4300 0.0000 132.6300 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279364 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279364 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[5]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 213.0210 155.1430 213.2210 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 213.0210 155.1430 213.2210 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 213.0210 155.1430 213.2210 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 213.0210 155.1430 213.2210 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 213.0210 155.1430 213.2210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.23524 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23524 LAYER M3 ;
    ANTENNAMAXAREACAR 22.98153 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 27.12209 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 31.26238 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[3]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 17.3160 155.1430 17.5160 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 17.3160 155.1430 17.5160 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 17.3160 155.1430 17.5160 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 17.3160 155.1430 17.5160 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 17.3160 155.1430 17.5160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.3739 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3739 LAYER M4 ;
    ANTENNAMAXAREACAR 16.1776 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 20.60928 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 9.8210 155.1430 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 9.8210 155.1430 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 9.8210 155.1430 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 9.8210 155.1430 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 9.8210 155.1430 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.64074 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.64074 LAYER M2 ;
    ANTENNAMAXAREACAR 12.26859 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 13.30542 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.34219 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.37889 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.9430 210.4120 155.1430 210.6120 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.9430 210.4120 155.1430 210.6120 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.9430 210.4120 155.1430 210.6120 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.9430 210.4120 155.1430 210.6120 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.9430 210.4120 155.1430 210.6120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.1830 0.0000 109.3830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.1830 0.0000 109.3830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.1830 0.0000 109.3830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.1830 0.0000 109.3830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.1830 0.0000 109.3830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[29]
  OBS
    LAYER M2 ;
      RECT 0.0000 255.3990 154.2490 261.5300 ;
      RECT 0.0000 229.9720 155.1430 255.3990 ;
      RECT 0.0000 228.3720 154.2430 229.9720 ;
      RECT 154.2430 211.3120 155.1430 212.3210 ;
      RECT 153.6420 258.1600 155.1430 259.9300 ;
      RECT 0.0000 221.4250 155.1430 228.3720 ;
      RECT 0.0000 219.0960 154.2430 221.4250 ;
      RECT 0.0000 213.9210 155.1430 219.0960 ;
      RECT 0.0000 209.7120 154.2430 213.9210 ;
      RECT 0.0000 203.8860 155.1430 209.7120 ;
      RECT 0.0000 201.6650 154.2430 203.8860 ;
      RECT 0.0000 51.8100 155.1430 201.6650 ;
      RECT 0.0000 50.2100 154.2430 51.8100 ;
      RECT 0.0000 18.2160 155.1430 50.2100 ;
      RECT 0.0000 16.1340 154.2430 18.2160 ;
      RECT 0.0000 10.7210 155.1430 16.1340 ;
      RECT 0.0000 9.1210 154.2430 10.7210 ;
      RECT 0.0000 0.9000 155.1430 9.1210 ;
      RECT 0.0000 0.0000 66.7750 0.9000 ;
      RECT 134.0390 0.0000 155.1430 9.1210 ;
      RECT 134.0390 0.0000 155.1430 0.9000 ;
      RECT 0.0000 261.5300 155.1430 268.1970 ;
      RECT 0.0000 229.9720 154.2490 268.1970 ;
      RECT 0.0000 0.0000 66.7750 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
    LAYER M1 ;
      RECT 154.3430 211.2120 155.1430 212.4210 ;
      RECT 153.6420 258.0600 155.1430 260.0300 ;
      RECT 0.0000 221.3250 155.1430 228.4720 ;
      RECT 0.0000 219.1960 154.3430 221.3250 ;
      RECT 0.0000 213.8210 155.1430 219.1960 ;
      RECT 0.0000 209.8120 154.3430 213.8210 ;
      RECT 0.0000 203.7860 155.1430 209.8120 ;
      RECT 0.0000 201.7650 154.3430 203.7860 ;
      RECT 0.0000 51.7100 155.1430 201.7650 ;
      RECT 0.0000 50.3100 154.3430 51.7100 ;
      RECT 0.0000 18.1160 155.1430 50.3100 ;
      RECT 0.0000 16.2340 154.3430 18.1160 ;
      RECT 0.0000 10.6210 155.1430 16.2340 ;
      RECT 0.0000 9.2210 154.3430 10.6210 ;
      RECT 0.0000 0.8000 155.1430 9.2210 ;
      RECT 0.0000 0.0000 66.8750 0.8000 ;
      RECT 133.9390 0.0000 155.1430 9.2210 ;
      RECT 133.9390 0.0000 155.1430 0.8000 ;
      RECT 0.0000 261.4300 155.1430 268.1970 ;
      RECT 0.0000 229.8720 154.3490 268.1970 ;
      RECT 0.0000 0.0000 66.8750 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 0.8000 154.3430 268.1970 ;
      RECT 0.0000 255.4990 154.3490 261.4300 ;
      RECT 0.0000 229.8720 155.1430 255.4990 ;
      RECT 0.0000 228.4720 154.3430 229.8720 ;
    LAYER PO ;
      RECT 0.0000 0.0000 155.1430 268.1970 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 155.1430 268.1970 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 155.1430 268.1970 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 155.1430 268.1970 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 155.1430 268.1970 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 155.1430 268.1970 ;
    LAYER M5 ;
      RECT 154.5580 267.1970 155.1430 268.1970 ;
      RECT 153.6420 258.1600 155.1430 259.9300 ;
      RECT 154.2430 211.3120 155.1430 212.3210 ;
      RECT 0.0000 221.4250 155.1430 228.3720 ;
      RECT 0.0000 219.0960 154.2430 221.4250 ;
      RECT 0.0000 213.9210 155.1430 219.0960 ;
      RECT 0.0000 209.7120 154.2430 213.9210 ;
      RECT 0.0000 203.8860 155.1430 209.7120 ;
      RECT 0.0000 201.6650 154.2430 203.8860 ;
      RECT 0.0000 51.8100 155.1430 201.6650 ;
      RECT 0.0000 50.2100 154.2430 51.8100 ;
      RECT 0.0000 18.2160 155.1430 50.2100 ;
      RECT 0.0000 16.1340 154.2430 18.2160 ;
      RECT 0.0000 10.7210 155.1430 16.1340 ;
      RECT 0.0000 9.1210 154.2430 10.7210 ;
      RECT 0.0000 0.9000 155.1430 9.1210 ;
      RECT 0.0000 0.0000 66.7750 0.9000 ;
      RECT 134.0390 0.0000 155.1430 9.1210 ;
      RECT 134.0390 0.0000 155.1430 0.9000 ;
      RECT 0.0000 261.5300 155.1430 267.1970 ;
      RECT 0.0000 229.9720 154.2490 267.1970 ;
      RECT 0.0000 0.0000 66.7750 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 0.9000 154.2430 267.1970 ;
      RECT 0.0000 255.3990 154.2490 261.5300 ;
      RECT 0.0000 229.9720 155.1430 255.3990 ;
      RECT 0.0000 228.3720 154.2430 229.9720 ;
    LAYER M4 ;
      RECT 154.2430 211.3120 155.1430 212.3210 ;
      RECT 153.6420 258.1600 155.1430 259.9300 ;
      RECT 0.0000 221.4250 155.1430 228.3720 ;
      RECT 0.0000 219.0960 154.2430 221.4250 ;
      RECT 0.0000 213.9210 155.1430 219.0960 ;
      RECT 0.0000 209.7120 154.2430 213.9210 ;
      RECT 0.0000 203.8860 155.1430 209.7120 ;
      RECT 0.0000 201.6650 154.2430 203.8860 ;
      RECT 0.0000 51.8100 155.1430 201.6650 ;
      RECT 0.0000 50.2100 154.2430 51.8100 ;
      RECT 0.0000 18.2160 155.1430 50.2100 ;
      RECT 0.0000 16.1340 154.2430 18.2160 ;
      RECT 0.0000 10.7210 155.1430 16.1340 ;
      RECT 0.0000 9.1210 154.2430 10.7210 ;
      RECT 0.0000 0.9000 155.1430 9.1210 ;
      RECT 0.0000 0.0000 66.7750 0.9000 ;
      RECT 134.0390 0.0000 155.1430 9.1210 ;
      RECT 134.0390 0.0000 155.1430 0.9000 ;
      RECT 0.0000 261.5300 155.1430 268.1970 ;
      RECT 0.0000 229.9720 154.2490 268.1970 ;
      RECT 0.0000 0.0000 66.7750 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 255.3990 154.2490 261.5300 ;
      RECT 0.0000 229.9720 155.1430 255.3990 ;
      RECT 0.0000 228.3720 154.2430 229.9720 ;
    LAYER M3 ;
      RECT 154.2430 211.3120 155.1430 212.3210 ;
      RECT 153.6420 258.1600 155.1430 259.9300 ;
      RECT 0.0000 221.4250 155.1430 228.3720 ;
      RECT 0.0000 219.0960 154.2430 221.4250 ;
      RECT 0.0000 213.9210 155.1430 219.0960 ;
      RECT 0.0000 209.7120 154.2430 213.9210 ;
      RECT 0.0000 203.8860 155.1430 209.7120 ;
      RECT 0.0000 201.6650 154.2430 203.8860 ;
      RECT 0.0000 51.8100 155.1430 201.6650 ;
      RECT 0.0000 50.2100 154.2430 51.8100 ;
      RECT 0.0000 18.2160 155.1430 50.2100 ;
      RECT 0.0000 16.1340 154.2430 18.2160 ;
      RECT 0.0000 10.7210 155.1430 16.1340 ;
      RECT 0.0000 9.1210 154.2430 10.7210 ;
      RECT 0.0000 0.9000 155.1430 9.1210 ;
      RECT 0.0000 0.0000 66.7750 0.9000 ;
      RECT 134.0390 0.0000 155.1430 9.1210 ;
      RECT 134.0390 0.0000 155.1430 0.9000 ;
      RECT 0.0000 261.5300 155.1430 268.1970 ;
      RECT 0.0000 229.9720 154.2490 268.1970 ;
      RECT 0.0000 0.0000 66.7750 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 0.9000 154.2430 268.1970 ;
      RECT 0.0000 255.3990 154.2490 261.5300 ;
      RECT 0.0000 229.9720 155.1430 255.3990 ;
      RECT 0.0000 228.3720 154.2430 229.9720 ;
  END
END SRAMLP1RW256x48

MACRO SRAMLP1RW256x128
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 372.879 BY 309.253 ;
  SYMMETRY X Y R90 ;

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 177.3690 0.0000 177.5690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.3690 0.0000 177.5690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.3690 0.0000 177.5690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 177.3690 0.0000 177.5690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 177.3690 0.0000 177.5690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[0]

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 358.2390 308.9530 358.5380 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 359.1390 308.9530 359.4390 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 360.0380 308.9530 360.3370 309.2530 ;
    END
  END VDDL

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 179.4200 0.0000 179.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.4200 0.0000 179.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.4200 0.0000 179.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 179.4200 0.0000 179.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 179.4200 0.0000 179.6200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 201.9930 0.0000 202.1930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 201.9930 0.0000 202.1930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 201.9930 0.0000 202.1930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 201.9930 0.0000 202.1930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 201.9930 0.0000 202.1930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[18]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.2040 0.0000 197.4040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.2040 0.0000 197.4040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.2040 0.0000 197.4040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.2040 0.0000 197.4040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.2040 0.0000 197.4040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 196.5210 0.0000 196.7210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 196.5210 0.0000 196.7210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 196.5210 0.0000 196.7210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 196.5210 0.0000 196.7210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 196.5210 0.0000 196.7210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[14]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 195.8360 0.0000 196.0360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 195.8360 0.0000 196.0360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 195.8360 0.0000 196.0360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 195.8360 0.0000 196.0360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 195.8360 0.0000 196.0360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 198.5720 0.0000 198.7720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 198.5720 0.0000 198.7720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 198.5720 0.0000 198.7720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 198.5720 0.0000 198.7720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 198.5720 0.0000 198.7720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.8890 0.0000 198.0890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.8890 0.0000 198.0890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.8890 0.0000 198.0890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.8890 0.0000 198.0890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.8890 0.0000 198.0890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[15]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 199.2570 0.0000 199.4570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 199.2570 0.0000 199.4570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 199.2570 0.0000 199.4570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 199.2570 0.0000 199.4570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 199.2570 0.0000 199.4570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[16]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 199.9400 0.0000 200.1400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 199.9400 0.0000 200.1400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 199.9400 0.0000 200.1400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 199.9400 0.0000 200.1400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 199.9400 0.0000 200.1400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 191.7320 0.0000 191.9320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 191.7320 0.0000 191.9320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 191.7320 0.0000 191.9320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 191.7320 0.0000 191.9320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 191.7320 0.0000 191.9320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 192.4170 0.0000 192.6170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 192.4170 0.0000 192.6170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 192.4170 0.0000 192.6170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 192.4170 0.0000 192.6170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 192.4170 0.0000 192.6170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[11]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 194.4680 0.0000 194.6680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 194.4680 0.0000 194.6680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 194.4680 0.0000 194.6680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 194.4680 0.0000 194.6680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 194.4680 0.0000 194.6680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 195.1530 0.0000 195.3530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 195.1530 0.0000 195.3530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 195.1530 0.0000 195.3530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 195.1530 0.0000 195.3530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 195.1530 0.0000 195.3530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[13]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 193.1000 0.0000 193.3000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 193.1000 0.0000 193.3000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 193.1000 0.0000 193.3000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 193.1000 0.0000 193.3000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 193.1000 0.0000 193.3000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 193.7850 0.0000 193.9850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 193.7850 0.0000 193.9850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 193.7850 0.0000 193.9850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 193.7850 0.0000 193.9850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 193.7850 0.0000 193.9850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[12]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 186.9450 0.0000 187.1450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.9450 0.0000 187.1450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.9450 0.0000 187.1450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 186.9450 0.0000 187.1450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 186.9450 0.0000 187.1450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[7]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 187.6280 0.0000 187.8280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 187.6280 0.0000 187.8280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 187.6280 0.0000 187.8280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 187.6280 0.0000 187.8280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 187.6280 0.0000 187.8280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 188.9960 0.0000 189.1960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 188.9960 0.0000 189.1960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 188.9960 0.0000 189.1960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 188.9960 0.0000 189.1960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 188.9960 0.0000 189.1960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 188.3130 0.0000 188.5130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 188.3130 0.0000 188.5130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 188.3130 0.0000 188.5130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 188.3130 0.0000 188.5130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 188.3130 0.0000 188.5130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[8]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 190.3640 0.0000 190.5640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.3640 0.0000 190.5640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.3640 0.0000 190.5640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 190.3640 0.0000 190.5640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 190.3640 0.0000 190.5640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 209.5160 0.0000 209.7160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 209.5160 0.0000 209.7160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 209.5160 0.0000 209.7160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 209.5160 0.0000 209.7160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 209.5160 0.0000 209.7160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 210.2010 0.0000 210.4010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 210.2010 0.0000 210.4010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 210.2010 0.0000 210.4010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 210.2010 0.0000 210.4010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 210.2010 0.0000 210.4010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[24]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 210.8840 0.0000 211.0840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 210.8840 0.0000 211.0840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 210.8840 0.0000 211.0840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 210.8840 0.0000 211.0840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 210.8840 0.0000 211.0840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 213.6200 0.0000 213.8200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 213.6200 0.0000 213.8200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 213.6200 0.0000 213.8200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 213.6200 0.0000 213.8200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 213.6200 0.0000 213.8200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 212.9370 0.0000 213.1370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.9370 0.0000 213.1370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.9370 0.0000 213.1370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 212.9370 0.0000 213.1370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 212.9370 0.0000 213.1370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[26]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 211.5690 0.0000 211.7690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.5690 0.0000 211.7690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.5690 0.0000 211.7690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 211.5690 0.0000 211.7690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 211.5690 0.0000 211.7690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[25]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 212.2520 0.0000 212.4520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.2520 0.0000 212.4520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.2520 0.0000 212.4520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 212.2520 0.0000 212.4520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 212.2520 0.0000 212.4520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 204.7290 0.0000 204.9290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.7290 0.0000 204.9290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.7290 0.0000 204.9290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 204.7290 0.0000 204.9290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 204.7290 0.0000 204.9290 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[20]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 205.4120 0.0000 205.6120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.4120 0.0000 205.6120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.4120 0.0000 205.6120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 205.4120 0.0000 205.6120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 205.4120 0.0000 205.6120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 206.0970 0.0000 206.2970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 206.0970 0.0000 206.2970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 206.0970 0.0000 206.2970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 206.0970 0.0000 206.2970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 206.0970 0.0000 206.2970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[21]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 207.4650 0.0000 207.6650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 207.4650 0.0000 207.6650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 207.4650 0.0000 207.6650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 207.4650 0.0000 207.6650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 207.4650 0.0000 207.6650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[22]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 208.1480 0.0000 208.3480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 208.1480 0.0000 208.3480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 208.1480 0.0000 208.3480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 208.1480 0.0000 208.3480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 208.1480 0.0000 208.3480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 206.7800 0.0000 206.9800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 206.7800 0.0000 206.9800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 206.7800 0.0000 206.9800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 206.7800 0.0000 206.9800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 206.7800 0.0000 206.9800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 201.3080 0.0000 201.5080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 201.3080 0.0000 201.5080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 201.3080 0.0000 201.5080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 201.3080 0.0000 201.5080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 201.3080 0.0000 201.5080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 200.6250 0.0000 200.8250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 200.6250 0.0000 200.8250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 200.6250 0.0000 200.8250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 200.6250 0.0000 200.8250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 200.6250 0.0000 200.8250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[17]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 204.0440 0.0000 204.2440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.0440 0.0000 204.2440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.0440 0.0000 204.2440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 204.0440 0.0000 204.2440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 204.0440 0.0000 204.2440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 202.6760 0.0000 202.8760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 202.6760 0.0000 202.8760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 202.6760 0.0000 202.8760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 202.6760 0.0000 202.8760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 202.6760 0.0000 202.8760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 203.3610 0.0000 203.5610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.3610 0.0000 203.5610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.3610 0.0000 203.5610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 203.3610 0.0000 203.5610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 203.3610 0.0000 203.5610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[19]

  PIN O[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 244.4010 0.0000 244.6010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 244.4010 0.0000 244.6010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 244.4010 0.0000 244.6010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 244.4010 0.0000 244.6010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 244.4010 0.0000 244.6010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[49]

  PIN I[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 243.7160 0.0000 243.9160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 243.7160 0.0000 243.9160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 243.7160 0.0000 243.9160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 243.7160 0.0000 243.9160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 243.7160 0.0000 243.9160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[49]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 9.8200 372.8790 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 9.8200 372.8790 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 9.8200 372.8790 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 9.8200 372.8790 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 9.8200 372.8790 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 240.2970 0.0000 240.4970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 240.2970 0.0000 240.4970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 240.2970 0.0000 240.4970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 240.2970 0.0000 240.4970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 240.2970 0.0000 240.4970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[46]

  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 239.6120 0.0000 239.8120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 239.6120 0.0000 239.8120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 239.6120 0.0000 239.8120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 239.6120 0.0000 239.8120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 239.6120 0.0000 239.8120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[46]

  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 240.9800 0.0010 241.1800 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 240.9800 0.0010 241.1800 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 240.9800 0.0000 241.1800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 240.9800 0.0000 241.1800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 240.9800 0.0000 241.1800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[47]

  PIN O[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 263.5530 0.0000 263.7530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 263.5530 0.0000 263.7530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 263.5530 0.0000 263.7530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 263.5530 0.0000 263.7530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 263.5530 0.0000 263.7530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[63]

  PIN I[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 262.8680 0.0000 263.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 262.8680 0.0000 263.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 262.8680 0.0000 263.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 262.8680 0.0000 263.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 262.8680 0.0000 263.0680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[63]

  PIN O[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 262.1850 0.0000 262.3850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 262.1850 0.0000 262.3850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 262.1850 0.0000 262.3850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 262.1850 0.0000 262.3850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 262.1850 0.0000 262.3850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[62]

  PIN I[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 261.5000 0.0000 261.7000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 261.5000 0.0000 261.7000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 261.5000 0.0000 261.7000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 261.5000 0.0000 261.7000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 261.5000 0.0000 261.7000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[62]

  PIN O[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 264.9210 0.0000 265.1210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 264.9210 0.0000 265.1210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 264.9210 0.0000 265.1210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 264.9210 0.0000 265.1210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 264.9210 0.0000 265.1210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[64]

  PIN I[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 264.2360 0.0000 264.4360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 264.2360 0.0000 264.4360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 264.2360 0.0000 264.4360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 264.2360 0.0000 264.4360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 264.2360 0.0000 264.4360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[64]

  PIN O[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 256.7130 0.0000 256.9130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 256.7130 0.0000 256.9130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 256.7130 0.0000 256.9130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 256.7130 0.0000 256.9130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 256.7130 0.0000 256.9130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[58]

  PIN I[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 256.0280 0.0000 256.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 256.0280 0.0000 256.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 256.0280 0.0000 256.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 256.0280 0.0000 256.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 256.0280 0.0000 256.2280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[58]

  PIN I[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 258.7640 0.0000 258.9640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 258.7640 0.0000 258.9640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 258.7640 0.0000 258.9640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 258.7640 0.0000 258.9640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 258.7640 0.0000 258.9640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[60]

  PIN O[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 260.8170 0.0000 261.0170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.8170 0.0000 261.0170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.8170 0.0000 261.0170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 260.8170 0.0000 261.0170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 260.8170 0.0000 261.0170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[61]

  PIN I[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 257.3960 0.0000 257.5960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 257.3960 0.0000 257.5960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 257.3960 0.0000 257.5960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 257.3960 0.0000 257.5960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 257.3960 0.0000 257.5960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[59]

  PIN O[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 258.0810 0.0000 258.2810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 258.0810 0.0000 258.2810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 258.0810 0.0000 258.2810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 258.0810 0.0000 258.2810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 258.0810 0.0000 258.2810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[59]

  PIN I[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 260.1320 0.0000 260.3320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.1320 0.0000 260.3320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.1320 0.0000 260.3320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 260.1320 0.0000 260.3320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 260.1320 0.0000 260.3320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[61]

  PIN O[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 259.4490 0.0000 259.6490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 259.4490 0.0000 259.6490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 259.4490 0.0000 259.6490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 259.4490 0.0000 259.6490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 259.4490 0.0000 259.6490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[60]

  PIN O[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 255.3450 0.0000 255.5450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.3450 0.0000 255.5450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.3450 0.0000 255.5450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 255.3450 0.0000 255.5450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 255.3450 0.0000 255.5450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[57]

  PIN O[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 253.9770 0.0000 254.1770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 253.9770 0.0000 254.1770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 253.9770 0.0000 254.1770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 253.9770 0.0000 254.1770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 253.9770 0.0000 254.1770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[56]

  PIN I[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 253.2920 0.0000 253.4920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 253.2920 0.0000 253.4920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 253.2920 0.0000 253.4920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 253.2920 0.0000 253.4920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 253.2920 0.0000 253.4920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[56]

  PIN I[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 254.6600 0.0000 254.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 254.6600 0.0000 254.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 254.6600 0.0000 254.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 254.6600 0.0000 254.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 254.6600 0.0000 254.8600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[57]

  PIN I[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 276.5480 0.0000 276.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 276.5480 0.0000 276.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 276.5480 0.0000 276.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 276.5480 0.0000 276.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 276.5480 0.0000 276.7480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[73]

  PIN O[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 277.2330 0.0000 277.4330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 277.2330 0.0000 277.4330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 277.2330 0.0000 277.4330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 277.2330 0.0000 277.4330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 277.2330 0.0000 277.4330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[73]

  PIN O[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 278.6010 0.0000 278.8010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.6010 0.0000 278.8010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.6010 0.0000 278.8010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 278.6010 0.0000 278.8010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 278.6010 0.0000 278.8010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[74]

  PIN I[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 277.9160 0.0000 278.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 277.9160 0.0000 278.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 277.9160 0.0000 278.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 277.9160 0.0000 278.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 277.9160 0.0000 278.1160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[74]

  PIN I[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 275.1800 0.0000 275.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 275.1800 0.0000 275.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 275.1800 0.0000 275.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 275.1800 0.0000 275.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 275.1800 0.0000 275.3800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[72]

  PIN O[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 274.4970 0.0000 274.6970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 274.4970 0.0000 274.6970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 274.4970 0.0000 274.6970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 274.4970 0.0000 274.6970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 274.4970 0.0000 274.6970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[71]

  PIN I[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 273.8120 0.0000 274.0120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 273.8120 0.0000 274.0120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 273.8120 0.0000 274.0120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 273.8120 0.0000 274.0120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 273.8120 0.0000 274.0120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[71]

  PIN O[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 273.1290 0.0000 273.3290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 273.1290 0.0000 273.3290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 273.1290 0.0000 273.3290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 273.1290 0.0000 273.3290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 273.1290 0.0000 273.3290 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[70]

  PIN I[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 269.7080 0.0000 269.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 269.7080 0.0000 269.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 269.7080 0.0000 269.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 269.7080 0.0000 269.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 269.7080 0.0000 269.9080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[68]

  PIN I[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 272.4440 0.0000 272.6440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 272.4440 0.0000 272.6440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 272.4440 0.0000 272.6440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 272.4440 0.0000 272.6440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 272.4440 0.0000 272.6440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[70]

  PIN O[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 271.7610 0.0000 271.9610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 271.7610 0.0000 271.9610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 271.7610 0.0000 271.9610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 271.7610 0.0000 271.9610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 271.7610 0.0000 271.9610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[69]

  PIN I[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 271.0760 0.0000 271.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 271.0760 0.0000 271.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 271.0760 0.0000 271.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 271.0760 0.0000 271.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 271.0760 0.0000 271.2760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[69]

  PIN O[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 270.3930 0.0000 270.5930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 270.3930 0.0000 270.5930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 270.3930 0.0000 270.5930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 270.3930 0.0000 270.5930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 270.3930 0.0000 270.5930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[68]

  PIN O[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 266.2890 0.0000 266.4890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 266.2890 0.0000 266.4890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 266.2890 0.0000 266.4890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 266.2890 0.0000 266.4890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 266.2890 0.0000 266.4890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[65]

  PIN I[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 265.6040 0.0000 265.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 265.6040 0.0000 265.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 265.6040 0.0000 265.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 265.6040 0.0000 265.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 265.6040 0.0000 265.8040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[65]

  PIN I[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 266.9720 0.0000 267.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 266.9720 0.0000 267.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 266.9720 0.0000 267.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 266.9720 0.0000 267.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 266.9720 0.0000 267.1720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[66]

  PIN O[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 269.0250 0.0000 269.2250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 269.0250 0.0000 269.2250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 269.0250 0.0000 269.2250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 269.0250 0.0000 269.2250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 269.0250 0.0000 269.2250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[67]

  PIN I[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 268.3400 0.0000 268.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 268.3400 0.0000 268.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 268.3400 0.0000 268.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 268.3400 0.0000 268.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 268.3400 0.0000 268.5400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[67]

  PIN O[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 267.6570 0.0000 267.8570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 267.6570 0.0000 267.8570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 267.6570 0.0000 267.8570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 267.6570 0.0000 267.8570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 267.6570 0.0000 267.8570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[66]

  PIN I[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 242.3480 0.0000 242.5480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 242.3480 0.0000 242.5480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 242.3480 0.0000 242.5480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 242.3480 0.0000 242.5480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 242.3480 0.0000 242.5480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[48]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6850 287.8530 372.8790 288.0530 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6850 287.8530 372.8790 288.0530 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6850 287.8530 372.8790 288.0530 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6850 287.8530 372.8790 288.0530 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6850 287.8530 372.8790 288.0530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 351.7780 0.0000 351.9780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 351.7780 0.0000 351.9780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 351.7780 0.0000 351.9780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 351.7780 0.0000 351.9780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 351.7780 0.0000 351.9780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 94.1160 372.8790 94.3160 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 94.1160 372.8790 94.3160 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 94.1160 372.8790 94.3160 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 94.1160 372.8790 94.3160 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 94.1160 372.8790 94.3160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN O[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 288.1770 0.0000 288.3770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 288.1770 0.0000 288.3770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 288.1770 0.0000 288.3770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 288.1770 0.0000 288.3770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 288.1770 0.0000 288.3770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[81]

  PIN O[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 285.4410 0.0000 285.6410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 285.4410 0.0000 285.6410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 285.4410 0.0000 285.6410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 285.4410 0.0000 285.6410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 285.4410 0.0000 285.6410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[79]

  PIN I[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 287.4920 0.0000 287.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 287.4920 0.0000 287.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 287.4920 0.0000 287.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 287.4920 0.0000 287.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 287.4920 0.0000 287.6920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[81]

  PIN I[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 284.7560 0.0000 284.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 284.7560 0.0000 284.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 284.7560 0.0000 284.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 284.7560 0.0000 284.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 284.7560 0.0000 284.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[79]

  PIN I[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 286.1240 0.0000 286.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 286.1240 0.0000 286.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 286.1240 0.0000 286.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 286.1240 0.0000 286.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 286.1240 0.0000 286.3240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[80]

  PIN O[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 286.8090 0.0000 287.0090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 286.8090 0.0000 287.0090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 286.8090 0.0000 287.0090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 286.8090 0.0000 287.0090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 286.8090 0.0000 287.0090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[80]

  PIN O[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 282.7050 0.0000 282.9050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 282.7050 0.0000 282.9050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 282.7050 0.0000 282.9050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 282.7050 0.0000 282.9050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 282.7050 0.0000 282.9050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[77]

  PIN I[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 283.3880 0.0000 283.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 283.3880 0.0000 283.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 283.3880 0.0000 283.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 283.3880 0.0000 283.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 283.3880 0.0000 283.5880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[78]

  PIN O[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 284.0730 0.0000 284.2730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 284.0730 0.0000 284.2730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 284.0730 0.0000 284.2730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 284.0730 0.0000 284.2730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 284.0730 0.0000 284.2730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[78]

  PIN I[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 282.0200 0.0000 282.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 282.0200 0.0000 282.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 282.0200 0.0000 282.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 282.0200 0.0000 282.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 282.0200 0.0000 282.2200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[77]

  PIN I[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 279.2840 0.0000 279.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 279.2840 0.0000 279.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 279.2840 0.0000 279.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 279.2840 0.0000 279.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 279.2840 0.0000 279.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[75]

  PIN O[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 279.9690 0.0000 280.1690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 279.9690 0.0000 280.1690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 279.9690 0.0000 280.1690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 279.9690 0.0000 280.1690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 279.9690 0.0000 280.1690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[75]

  PIN I[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 280.6520 0.0000 280.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 280.6520 0.0000 280.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 280.6520 0.0000 280.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 280.6520 0.0000 280.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 280.6520 0.0000 280.8520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[76]

  PIN O[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 281.3370 0.0000 281.5370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 281.3370 0.0000 281.5370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 281.3370 0.0000 281.5370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 281.3370 0.0000 281.5370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 281.3370 0.0000 281.5370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[76]

  PIN O[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 275.8650 0.0000 276.0650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 275.8650 0.0000 276.0650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 275.8650 0.0000 276.0650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 275.8650 0.0000 276.0650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 275.8650 0.0000 276.0650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[72]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 189.6810 0.0000 189.8810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 189.6810 0.0000 189.8810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 189.6810 0.0000 189.8810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 189.6810 0.0000 189.8810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 189.6810 0.0000 189.8810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[9]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 191.0490 0.0000 191.2490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 191.0490 0.0000 191.2490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 191.0490 0.0000 191.2490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 191.0490 0.0000 191.2490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 191.0490 0.0000 191.2490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[10]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 183.5240 0.0000 183.7240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.5240 0.0000 183.7240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.5240 0.0000 183.7240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 183.5240 0.0000 183.7240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 183.5240 0.0000 183.7240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 184.2090 0.0000 184.4090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 184.2090 0.0000 184.4090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 184.2090 0.0000 184.4090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 184.2090 0.0000 184.4090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 184.2090 0.0000 184.4090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[5]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 182.8410 0.0000 183.0410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.8410 0.0000 183.0410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.8410 0.0000 183.0410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 182.8410 0.0000 183.0410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 182.8410 0.0000 183.0410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[4]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 184.8920 0.0000 185.0920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 184.8920 0.0000 185.0920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 184.8920 0.0000 185.0920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 184.8920 0.0000 185.0920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 184.8920 0.0000 185.0920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 185.5770 0.0000 185.7770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 185.5770 0.0000 185.7770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 185.5770 0.0000 185.7770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 185.5770 0.0000 185.7770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 185.5770 0.0000 185.7770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[6]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 186.2600 0.0000 186.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.2600 0.0000 186.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.2600 0.0000 186.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 186.2600 0.0000 186.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 186.2600 0.0000 186.4600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 178.7370 0.0000 178.9370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.7370 0.0000 178.9370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.7370 0.0000 178.9370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 178.7370 0.0000 178.9370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 178.7370 0.0000 178.9370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[1]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6850 288.1960 372.8790 288.3960 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6850 288.1960 372.8790 288.3960 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6850 288.1960 372.8790 288.3960 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6850 288.1960 372.8790 288.3960 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6850 288.1960 372.8790 288.3960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 180.7880 0.0000 180.9880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 180.7880 0.0000 180.9880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 180.7880 0.0000 180.9880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 180.7880 0.0000 180.9880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 180.7880 0.0000 180.9880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 181.4730 0.0000 181.6730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 181.4730 0.0000 181.6730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 181.4730 0.0000 181.6730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 181.4730 0.0000 181.6730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 181.4730 0.0000 181.6730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[3]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 182.1560 0.0000 182.3560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.1560 0.0000 182.3560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.1560 0.0000 182.3560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 182.1560 0.0000 182.3560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 182.1560 0.0000 182.3560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 180.1050 0.0000 180.3050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 180.1050 0.0000 180.3050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 180.1050 0.0000 180.3050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 180.1050 0.0000 180.3050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 180.1050 0.0000 180.3050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[2]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 178.0520 0.0010 178.2520 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.0520 0.0010 178.2520 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.0520 0.0000 178.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 178.0520 0.0000 178.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 178.0520 0.0000 178.2520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 176.6840 0.0000 176.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.6840 0.0000 176.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.6840 0.0000 176.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 176.6840 0.0000 176.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 176.6840 0.0000 176.8840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 350.4200 0.0000 350.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 350.4200 0.0000 350.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 350.4200 0.0000 350.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 350.4200 0.0000 350.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 350.4200 0.0000 350.6200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[127]

  PIN O[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 351.1050 0.0000 351.3050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 351.1050 0.0000 351.3050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 351.1050 0.0000 351.3050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 351.1050 0.0000 351.3050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 351.1050 0.0000 351.3050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[127]

  PIN O[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 347.0010 0.0000 347.2010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 347.0010 0.0000 347.2010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 347.0010 0.0000 347.2010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 347.0010 0.0000 347.2010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 347.0010 0.0000 347.2010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[124]

  PIN I[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 349.0520 0.0000 349.2520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 349.0520 0.0000 349.2520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 349.0520 0.0000 349.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 349.0520 0.0000 349.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 349.0520 0.0000 349.2520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[126]

  PIN I[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 346.3160 0.0000 346.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 346.3160 0.0000 346.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 346.3160 0.0000 346.5160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 346.3160 0.0000 346.5160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 346.3160 0.0000 346.5160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[124]

  PIN I[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 347.6840 0.0000 347.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 347.6840 0.0000 347.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 347.6840 0.0000 347.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 347.6840 0.0000 347.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 347.6840 0.0000 347.8840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[125]

  PIN O[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 345.6330 0.0000 345.8330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 345.6330 0.0000 345.8330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 345.6330 0.0000 345.8330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 345.6330 0.0000 345.8330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 345.6330 0.0000 345.8330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[123]

  PIN O[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 348.3690 0.0000 348.5690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 348.3690 0.0000 348.5690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 348.3690 0.0000 348.5690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 348.3690 0.0000 348.5690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 348.3690 0.0000 348.5690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[125]

  PIN O[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 342.8970 0.0000 343.0970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 342.8970 0.0000 343.0970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 342.8970 0.0000 343.0970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 342.8970 0.0000 343.0970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 342.8970 0.0000 343.0970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[121]

  PIN I[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 344.9480 0.0000 345.1480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 344.9480 0.0000 345.1480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 344.9480 0.0000 345.1480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 344.9480 0.0000 345.1480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 344.9480 0.0000 345.1480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[123]

  PIN I[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 342.2120 0.0000 342.4120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 342.2120 0.0000 342.4120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 342.2120 0.0000 342.4120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 342.2120 0.0000 342.4120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 342.2120 0.0000 342.4120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[121]

  PIN O[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 341.5290 0.0000 341.7290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 341.5290 0.0000 341.7290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 341.5290 0.0000 341.7290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 341.5290 0.0000 341.7290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 341.5290 0.0000 341.7290 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[120]

  PIN O[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 344.2650 0.0000 344.4650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 344.2650 0.0000 344.4650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 344.2650 0.0000 344.4650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 344.2650 0.0000 344.4650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 344.2650 0.0000 344.4650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[122]

  PIN I[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 343.5800 0.0000 343.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 343.5800 0.0000 343.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 343.5800 0.0000 343.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 343.5800 0.0000 343.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 343.5800 0.0000 343.7800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[122]

  PIN O[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 338.7930 0.0000 338.9930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 338.7930 0.0000 338.9930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 338.7930 0.0000 338.9930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 338.7930 0.0000 338.9930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 338.7930 0.0000 338.9930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[118]

  PIN I[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 338.1080 0.0000 338.3080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 338.1080 0.0000 338.3080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 338.1080 0.0000 338.3080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 338.1080 0.0000 338.3080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 338.1080 0.0000 338.3080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[118]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 264.8010 372.8790 265.0010 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 264.8010 372.8790 265.0010 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 264.8010 372.8790 265.0010 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 264.8010 372.8790 265.0010 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 264.8010 372.8790 265.0010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 245.5750 372.8790 245.7750 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 245.5750 372.8790 245.7750 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 245.5750 372.8790 245.7750 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 245.5750 372.8790 245.7750 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 245.5750 372.8790 245.7750 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6850 291.4480 372.8790 291.6480 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6850 291.4480 372.8790 291.6480 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6850 291.4480 372.8790 291.6480 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6850 291.4480 372.8790 291.6480 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6850 291.4480 372.8790 291.6480 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 219.0920 0.0000 219.2920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.0920 0.0000 219.2920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.0920 0.0000 219.2920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 219.0920 0.0000 219.2920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 219.0920 0.0000 219.2920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 218.4090 0.0000 218.6090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 218.4090 0.0000 218.6090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 218.4090 0.0000 218.6090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 218.4090 0.0000 218.6090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 218.4090 0.0000 218.6090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[30]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 208.8330 0.0000 209.0330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 208.8330 0.0000 209.0330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 208.8330 0.0000 209.0330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 208.8330 0.0000 209.0330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 208.8330 0.0000 209.0330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[23]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 247.1650 372.8790 247.3650 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 247.1650 372.8790 247.3650 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 247.1650 372.8790 247.3650 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 247.1650 372.8790 247.3650 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 247.1650 372.8790 247.3650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 254.3910 372.8790 254.5910 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 254.3910 372.8790 254.5910 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 254.3910 372.8790 254.5910 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 254.3910 372.8790 254.5910 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 254.3910 372.8790 254.5910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 255.9810 372.8790 256.1810 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 255.9810 372.8790 256.1810 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 255.9810 372.8790 256.1810 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 255.9810 372.8790 256.1810 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 255.9810 372.8790 256.1810 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 263.2110 372.8790 263.4110 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 263.2110 372.8790 263.4110 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 263.2110 372.8790 263.4110 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 263.2110 372.8790 263.4110 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 263.2110 372.8790 263.4110 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 272.0310 372.8790 272.2310 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 272.0310 372.8790 272.2310 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 272.0310 372.8790 272.2310 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 272.0310 372.8790 272.2310 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 272.0310 372.8790 272.2310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 369.0380 308.9530 369.3370 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 370.8370 308.9530 371.1360 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 369.9380 308.9530 370.2380 309.2530 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.0900 308.9530 4.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2900 308.9530 2.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.1910 308.9530 3.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3900 308.9530 1.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.4910 308.9530 0.7920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.5900 308.9530 8.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.6900 308.9530 7.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8900 308.9530 6.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9900 308.9530 5.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.7910 308.9530 7.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.0890 308.9530 13.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1900 308.9530 12.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.2900 308.9530 11.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.4900 308.9530 9.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.9900 308.9530 14.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.3910 308.9530 10.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.6910 308.9530 16.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.7910 308.9530 16.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4900 308.9530 18.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.8890 308.9530 15.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.5910 308.9530 17.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.2900 308.9530 20.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.0910 308.9530 22.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.9900 308.9530 23.2890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.3900 308.9530 19.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.1900 308.9530 21.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.8910 308.9530 24.1920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.5910 308.9530 26.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.3910 308.9530 28.6920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.4900 308.9530 27.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.7900 308.9530 25.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.6900 308.9530 25.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.2900 308.9530 29.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.8910 308.9530 33.1920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.1900 308.9530 30.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.9900 308.9530 32.2890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.0910 308.9530 31.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.3900 308.9530 37.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.4900 308.9530 36.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.6900 308.9530 34.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.5910 308.9530 35.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.7900 308.9530 34.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.8900 308.9530 42.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.9900 308.9530 41.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.0900 308.9530 40.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.2900 308.9530 38.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.7910 308.9530 43.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.1910 308.9530 39.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.2890 308.9530 47.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.4890 308.9530 45.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.5900 308.9530 44.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.6900 308.9530 43.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.3900 308.9530 46.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.0910 308.9530 49.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.1910 308.9530 48.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.8900 308.9530 51.1910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.7900 308.9530 52.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.9910 308.9530 50.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.6900 308.9530 52.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.2910 308.9530 56.5920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.4910 308.9530 54.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.3900 308.9530 55.6890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.1900 308.9530 57.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.5900 308.9530 53.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.6900 308.9530 61.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.9910 308.9530 59.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.7910 308.9530 61.0920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.8900 308.9530 60.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.0900 308.9530 58.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.0900 308.9530 67.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.1900 308.9530 66.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.2910 308.9530 65.5920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.5900 308.9530 62.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.3900 308.9530 64.6890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.4910 308.9530 63.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.6900 308.9530 70.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.7900 308.9530 70.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.8900 308.9530 69.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.5910 308.9530 71.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.9910 308.9530 68.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.0900 308.9530 76.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.2900 308.9530 74.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.3900 308.9530 73.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.4900 308.9530 72.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.1910 308.9530 75.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.4910 308.9530 81.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.5910 308.9530 80.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.6890 308.9530 79.9890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.8890 308.9530 78.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.9900 308.9530 77.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.7900 308.9530 79.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.0900 308.9530 85.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.2900 308.9530 83.5910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.1900 308.9530 84.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.9900 308.9530 86.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.3910 308.9530 82.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.6910 308.9530 88.9920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.8910 308.9530 87.1910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.7900 308.9530 88.0890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.5900 308.9530 89.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.4900 308.9530 90.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.0900 308.9530 94.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.3910 308.9530 91.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.1910 308.9530 93.4920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.2900 308.9530 92.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.9900 308.9530 95.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.8910 308.9530 96.1910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.4900 308.9530 99.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.3910 308.9530 100.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.5900 308.9530 98.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.6910 308.9530 97.9920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.7900 308.9530 97.0890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.7900 308.9530 106.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.8900 308.9530 105.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.0900 308.9530 103.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.1900 308.9530 102.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.2900 308.9530 101.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.9910 308.9530 104.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.2890 308.9530 110.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.3900 308.9530 109.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.4900 308.9530 108.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.6900 308.9530 106.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.5910 308.9530 107.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.8910 308.9530 114.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.9910 308.9530 113.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.0890 308.9530 112.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.1900 308.9530 111.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.7910 308.9530 115.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.4900 308.9530 117.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.6900 308.9530 115.9910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.2910 308.9530 119.5910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.1900 308.9530 120.4890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.5900 308.9530 116.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.3900 308.9530 118.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.0910 308.9530 121.3920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.7910 308.9530 124.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.6900 308.9530 124.9890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.9900 308.9530 122.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.8900 308.9530 123.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.4900 308.9530 126.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.5910 308.9530 125.8920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.3900 308.9530 127.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.1900 308.9530 129.4890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.2910 308.9530 128.5910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.5900 308.9530 134.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.6900 308.9530 133.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.8900 308.9530 132.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.7910 308.9530 133.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.9900 308.9530 131.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.0910 308.9530 130.3920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.0900 308.9530 139.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.1900 308.9530 138.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.2900 308.9530 137.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.4900 308.9530 135.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.3910 308.9530 136.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.6890 308.9530 142.9890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.7900 308.9530 142.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.8900 308.9530 141.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.5900 308.9530 143.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.9910 308.9530 140.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.2910 308.9530 146.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.3910 308.9530 145.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.0900 308.9530 148.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.4890 308.9530 144.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.9900 308.9530 149.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.1910 308.9530 147.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.8900 308.9530 150.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.6910 308.9530 151.9910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.5900 308.9530 152.8890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.4910 308.9530 153.7920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.7900 308.9530 151.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.8900 308.9530 159.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.1910 308.9530 156.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.9910 308.9530 158.2920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.0900 308.9530 157.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.3900 308.9530 154.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.2900 308.9530 155.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 163.3900 308.9530 163.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.4910 308.9530 162.7920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.7900 308.9530 160.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.5900 308.9530 161.8890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.6910 308.9530 160.9910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.8900 308.9530 168.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.9900 308.9530 167.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.0900 308.9530 166.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.2900 308.9530 164.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.1910 308.9530 165.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.2900 308.9530 173.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.4900 308.9530 171.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.5900 308.9530 170.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.6900 308.9530 169.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.3910 308.9530 172.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.7910 308.9530 169.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.7910 308.9530 178.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.8890 308.9530 177.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.0890 308.9530 175.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 174.1900 308.9530 174.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.9900 308.9530 176.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.6910 308.9530 178.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.2900 308.9530 182.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.4900 308.9530 180.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.3900 308.9530 181.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.5910 308.9530 179.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.0910 308.9530 184.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.9900 308.9530 185.2890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.7900 308.9530 187.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 185.8910 308.9530 186.1920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.1900 308.9530 183.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 187.6900 308.9530 187.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.2900 308.9530 191.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.5910 308.9530 188.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.3910 308.9530 190.6920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.4900 308.9530 189.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.1900 308.9530 192.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.6900 308.9530 196.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.5910 308.9530 197.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 195.7900 308.9530 196.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.8910 308.9530 195.1920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.9900 308.9530 194.2890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.0910 308.9530 193.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 202.0900 308.9530 202.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 200.2900 308.9530 200.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 199.3900 308.9530 199.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 198.4900 308.9530 198.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 201.1910 308.9530 201.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 206.5900 308.9530 206.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.6900 308.9530 205.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.8900 308.9530 204.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 202.9900 308.9530 203.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.7910 308.9530 205.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.0910 308.9530 211.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 210.1910 308.9530 210.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 209.2890 308.9530 209.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.4890 308.9530 207.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 208.3900 308.9530 208.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.9910 308.9530 212.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 214.6900 308.9530 214.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.8900 308.9530 213.1910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.4910 308.9530 216.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 213.7900 308.9530 214.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.5900 308.9530 215.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.9910 308.9530 221.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 217.3900 308.9530 217.6890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.1900 308.9530 219.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 218.2910 308.9530 218.5920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.0900 308.9530 220.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 223.6900 308.9530 223.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.7910 308.9530 223.0920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 221.8900 308.9530 222.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 224.5900 308.9530 224.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.3900 308.9530 226.6890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 225.4910 308.9530 225.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.8900 308.9530 231.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 229.0900 308.9530 229.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 229.9910 308.9530 230.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.1900 308.9530 228.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 227.2910 308.9530 227.5920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 236.2900 308.9530 236.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 235.3900 308.9530 235.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.4900 308.9530 234.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 232.6900 308.9530 232.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 231.7900 308.9530 232.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.5910 308.9530 233.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 239.8890 308.9530 240.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 238.9900 308.9530 239.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 238.0900 308.9530 238.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 240.7900 308.9530 241.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 237.1910 308.9530 237.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 243.4910 308.9530 243.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 242.5910 308.9530 242.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 245.2900 308.9530 245.5910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.6890 308.9530 241.9890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 244.3910 308.9530 244.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 247.0900 308.9530 247.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.8910 308.9530 249.1910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 249.7900 308.9530 250.0890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 250.6910 308.9530 250.9920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 246.1900 308.9530 246.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 247.9900 308.9530 248.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 253.3910 308.9530 253.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.1910 308.9530 255.4920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 254.2900 308.9530 254.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 251.5900 308.9530 251.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 252.4900 308.9530 252.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 256.0900 308.9530 256.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 259.6910 308.9530 259.9920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 256.9900 308.9530 257.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 258.7900 308.9530 259.0890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 257.8910 308.9530 258.1910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 265.0900 308.9530 265.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 264.1900 308.9530 264.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 263.2900 308.9530 263.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 261.4900 308.9530 261.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 262.3910 308.9530 262.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.5900 308.9530 260.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 268.6900 308.9530 268.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 267.7900 308.9530 268.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 266.8900 308.9530 267.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 269.5910 308.9530 269.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 265.9910 308.9530 266.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 274.0890 308.9530 274.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 272.2890 308.9530 272.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 271.3900 308.9530 271.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 270.4900 308.9530 270.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 273.1900 308.9530 273.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 275.8910 308.9530 276.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 274.9910 308.9530 275.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 279.4900 308.9530 279.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 277.6900 308.9530 277.9910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.5900 308.9530 278.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 276.7910 308.9530 277.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 281.2910 308.9530 281.5910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 282.1900 308.9530 282.4890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 283.9900 308.9530 284.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 283.0910 308.9530 283.3920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 280.3900 308.9530 280.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 285.7910 308.9530 286.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 287.5910 308.9530 287.8920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 286.6900 308.9530 286.9890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 289.3900 308.9530 289.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 284.8900 308.9530 285.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 288.4900 308.9530 288.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 293.8900 308.9530 294.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 292.9900 308.9530 293.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 292.0910 308.9530 292.3920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 291.1900 308.9530 291.4890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 290.2910 308.9530 290.5910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 297.4900 308.9530 297.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 296.5900 308.9530 296.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 295.6900 308.9530 295.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 298.3910 308.9530 298.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 294.7910 308.9530 295.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 301.9910 308.9530 302.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 303.7900 308.9530 304.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 302.8900 308.9530 303.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 301.0900 308.9530 301.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 300.1900 308.9530 300.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 299.2900 308.9530 299.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 308.2910 308.9530 308.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 307.3910 308.9530 307.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 305.5900 308.9530 305.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 306.4890 308.9530 306.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 304.6890 308.9530 304.9890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 311.8900 308.9530 312.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.0900 308.9530 310.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.9900 308.9530 311.2910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 312.7900 308.9530 313.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 309.1910 308.9530 309.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 313.6910 308.9530 313.9910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 318.1910 308.9530 318.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 314.5900 308.9530 314.8890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 316.3900 308.9530 316.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 315.4910 308.9530 315.7920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 317.2900 308.9530 317.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 319.9910 308.9530 320.2920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 319.0900 308.9530 319.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 321.7900 308.9530 322.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 322.6910 308.9530 322.9910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 320.8900 308.9530 321.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 327.1910 308.9530 327.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 325.3900 308.9530 325.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 328.0900 308.9530 328.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 326.2900 308.9530 326.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 324.4910 308.9530 324.7920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 323.5900 308.9530 323.8890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 330.7910 308.9530 331.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 332.5900 308.9530 332.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 331.6900 308.9530 331.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 329.8900 308.9530 330.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 328.9900 308.9530 329.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 334.3910 308.9530 334.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 337.0890 308.9530 337.3890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 336.1900 308.9530 336.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 335.2900 308.9530 335.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 333.4900 308.9530 333.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 340.6910 308.9530 340.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 339.7910 308.9530 340.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 342.4900 308.9530 342.7910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 337.9900 308.9530 338.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 338.8890 308.9530 339.1890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 341.5910 308.9530 341.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 344.2900 308.9530 344.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 346.0910 308.9530 346.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 346.9900 308.9530 347.2890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 343.3900 308.9530 343.6910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 345.1900 308.9530 345.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 350.5910 308.9530 350.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 351.4900 308.9530 351.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 348.7900 308.9530 349.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 347.8910 308.9530 348.1920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 349.6900 308.9530 349.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 356.8910 308.9530 357.1920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 352.3910 308.9530 352.6920 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 354.1900 308.9530 354.4900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 355.9900 308.9530 356.2890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 355.0910 308.9530 355.3910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 353.2900 308.9530 353.5900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 359.5910 308.9530 359.8910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 357.7900 308.9530 358.0900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 361.3900 308.9530 361.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 360.4900 308.9530 360.7900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 358.6900 308.9530 358.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 363.1910 308.9530 363.4910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 365.8900 308.9530 366.1900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 364.9900 308.9530 365.2900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 364.0900 308.9530 364.3900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 367.6900 308.9530 367.9900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 368.5900 308.9530 368.8900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 369.4890 308.9530 369.7890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 371.2890 308.9530 371.5890 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 366.7910 308.9530 367.0910 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 370.3900 308.9530 370.6900 309.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 362.2900 308.9530 362.5900 309.2530 ;
    END
  END VSS

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 227.3000 0.0000 227.5000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 227.3000 0.0000 227.5000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 227.3000 0.0000 227.5000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 227.3000 0.0000 227.5000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 227.3000 0.0000 227.5000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[37]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 229.3530 0.0000 229.5530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 229.3530 0.0000 229.5530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 229.3530 0.0000 229.5530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 229.3530 0.0000 229.5530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 229.3530 0.0000 229.5530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[38]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 227.9850 0.0000 228.1850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 227.9850 0.0000 228.1850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 227.9850 0.0000 228.1850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 227.9850 0.0000 228.1850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 227.9850 0.0000 228.1850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[37]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 228.6680 0.0000 228.8680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.6680 0.0000 228.8680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.6680 0.0000 228.8680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 228.6680 0.0000 228.8680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 228.6680 0.0000 228.8680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 219.7770 0.0000 219.9770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.7770 0.0000 219.9770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.7770 0.0000 219.9770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 219.7770 0.0000 219.9770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 219.7770 0.0000 219.9770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[31]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 220.4600 0.0000 220.6600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 220.4600 0.0000 220.6600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 220.4600 0.0000 220.6600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 220.4600 0.0000 220.6600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 220.4600 0.0000 220.6600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 221.1450 0.0000 221.3450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 221.1450 0.0000 221.3450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 221.1450 0.0000 221.3450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 221.1450 0.0000 221.3450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 221.1450 0.0000 221.3450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[32]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 222.5130 0.0000 222.7130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 222.5130 0.0000 222.7130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 222.5130 0.0000 222.7130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 222.5130 0.0000 222.7130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 222.5130 0.0000 222.7130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[33]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 223.1960 0.0000 223.3960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 223.1960 0.0000 223.3960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 223.1960 0.0000 223.3960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 223.1960 0.0000 223.3960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 223.1960 0.0000 223.3960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 224.5640 0.0000 224.7640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 224.5640 0.0000 224.7640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 224.5640 0.0000 224.7640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 224.5640 0.0000 224.7640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 224.5640 0.0000 224.7640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 221.8280 0.0000 222.0280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 221.8280 0.0000 222.0280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 221.8280 0.0000 222.0280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 221.8280 0.0000 222.0280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 221.8280 0.0000 222.0280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 223.8810 0.0000 224.0810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 223.8810 0.0000 224.0810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 223.8810 0.0000 224.0810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 223.8810 0.0000 224.0810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 223.8810 0.0000 224.0810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[34]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 214.3050 0.0000 214.5050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 214.3050 0.0000 214.5050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 214.3050 0.0000 214.5050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 214.3050 0.0000 214.5050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 214.3050 0.0000 214.5050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[27]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 216.3560 0.0000 216.5560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 216.3560 0.0000 216.5560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 216.3560 0.0000 216.5560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 216.3560 0.0000 216.5560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 216.3560 0.0000 216.5560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 215.6730 0.0000 215.8730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.6730 0.0000 215.8730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.6730 0.0000 215.8730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 215.6730 0.0000 215.8730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 215.6730 0.0000 215.8730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[28]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 217.0410 0.0000 217.2410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 217.0410 0.0000 217.2410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 217.0410 0.0000 217.2410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 217.0410 0.0000 217.2410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 217.0410 0.0000 217.2410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[29]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 217.7240 0.0000 217.9240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 217.7240 0.0000 217.9240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 217.7240 0.0000 217.9240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 217.7240 0.0000 217.9240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 217.7240 0.0000 217.9240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 214.9880 0.0000 215.1880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 214.9880 0.0000 215.1880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 214.9880 0.0000 215.1880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 214.9880 0.0000 215.1880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 214.9880 0.0000 215.1880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 241.6650 0.0000 241.8650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.6650 0.0000 241.8650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.6650 0.0000 241.8650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 241.6650 0.0000 241.8650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 241.6650 0.0000 241.8650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[47]

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 237.5610 0.0000 237.7610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 237.5610 0.0000 237.7610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 237.5610 0.0000 237.7610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 237.5610 0.0000 237.7610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 237.5610 0.0000 237.7610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[44]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 234.8250 0.0000 235.0250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.8250 0.0000 235.0250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.8250 0.0000 235.0250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 234.8250 0.0000 235.0250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 234.8250 0.0000 235.0250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[42]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 235.5080 0.0000 235.7080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 235.5080 0.0000 235.7080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 235.5080 0.0000 235.7080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 235.5080 0.0000 235.7080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 235.5080 0.0000 235.7080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 236.1930 0.0000 236.3930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 236.1930 0.0000 236.3930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 236.1930 0.0000 236.3930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 236.1930 0.0000 236.3930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 236.1930 0.0000 236.3930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[43]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 236.8760 0.0000 237.0760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 236.8760 0.0000 237.0760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 236.8760 0.0000 237.0760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 236.8760 0.0000 237.0760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 236.8760 0.0000 237.0760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 238.2440 0.0000 238.4440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 238.2440 0.0000 238.4440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 238.2440 0.0000 238.4440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 238.2440 0.0000 238.4440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 238.2440 0.0000 238.4440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 238.9290 0.0000 239.1290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 238.9290 0.0000 239.1290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 238.9290 0.0000 239.1290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 238.9290 0.0000 239.1290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 238.9290 0.0000 239.1290 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[45]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 230.0360 0.0000 230.2360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.0360 0.0000 230.2360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.0360 0.0000 230.2360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 230.0360 0.0000 230.2360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 230.0360 0.0000 230.2360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[39]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 230.7210 0.0000 230.9210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.7210 0.0000 230.9210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.7210 0.0000 230.9210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 230.7210 0.0000 230.9210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 230.7210 0.0000 230.9210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[39]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 234.1400 0.0000 234.3400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.1400 0.0000 234.3400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.1400 0.0000 234.3400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 234.1400 0.0000 234.3400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 234.1400 0.0000 234.3400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[42]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 231.4040 0.0000 231.6040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 231.4040 0.0000 231.6040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 231.4040 0.0000 231.6040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 231.4040 0.0000 231.6040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 231.4040 0.0000 231.6040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[40]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 232.0890 0.0000 232.2890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 232.0890 0.0000 232.2890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 232.0890 0.0000 232.2890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 232.0890 0.0000 232.2890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 232.0890 0.0000 232.2890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[40]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 233.4570 0.0000 233.6570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.4570 0.0000 233.6570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.4570 0.0000 233.6570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 233.4570 0.0000 233.6570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 233.4570 0.0000 233.6570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[41]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 232.7720 0.0000 232.9720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 232.7720 0.0000 232.9720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 232.7720 0.0000 232.9720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 232.7720 0.0000 232.9720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 232.7720 0.0000 232.9720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[41]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 225.9320 0.0000 226.1320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 225.9320 0.0000 226.1320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 225.9320 0.0000 226.1320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 225.9320 0.0000 226.1320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 225.9320 0.0000 226.1320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 225.2490 0.0000 225.4490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 225.2490 0.0000 225.4490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 225.2490 0.0000 225.4490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 225.2490 0.0000 225.4490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 225.2490 0.0000 225.4490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[35]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 226.6170 0.0000 226.8170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.6170 0.0000 226.8170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.6170 0.0000 226.8170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 226.6170 0.0000 226.8170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 226.6170 0.0000 226.8170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[36]

  PIN O[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 252.6090 0.0000 252.8090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 252.6090 0.0000 252.8090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 252.6090 0.0000 252.8090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 252.6090 0.0000 252.8090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 252.6090 0.0000 252.8090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[55]

  PIN O[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 251.2410 0.0000 251.4410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 251.2410 0.0000 251.4410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 251.2410 0.0000 251.4410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 251.2410 0.0000 251.4410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 251.2410 0.0000 251.4410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[54]

  PIN I[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 251.9240 0.0000 252.1240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 251.9240 0.0000 252.1240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 251.9240 0.0000 252.1240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 251.9240 0.0000 252.1240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 251.9240 0.0000 252.1240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[55]

  PIN I[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 249.1880 0.0000 249.3880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 249.1880 0.0000 249.3880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 249.1880 0.0000 249.3880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 249.1880 0.0000 249.3880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 249.1880 0.0000 249.3880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[53]

  PIN O[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 248.5050 0.0000 248.7050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.5050 0.0000 248.7050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.5050 0.0000 248.7050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 248.5050 0.0000 248.7050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 248.5050 0.0000 248.7050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[52]

  PIN I[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 250.5560 0.0000 250.7560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 250.5560 0.0000 250.7560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 250.5560 0.0000 250.7560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 250.5560 0.0000 250.7560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 250.5560 0.0000 250.7560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[54]

  PIN O[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 249.8730 0.0000 250.0730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 249.8730 0.0000 250.0730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 249.8730 0.0000 250.0730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 249.8730 0.0000 250.0730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 249.8730 0.0000 250.0730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[53]

  PIN I[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 247.8200 0.0000 248.0200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 247.8200 0.0000 248.0200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 247.8200 0.0000 248.0200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 247.8200 0.0000 248.0200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 247.8200 0.0000 248.0200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[52]

  PIN O[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 247.1370 0.0000 247.3370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 247.1370 0.0000 247.3370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 247.1370 0.0000 247.3370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 247.1370 0.0000 247.3370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 247.1370 0.0000 247.3370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[51]

  PIN O[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 245.7690 0.0000 245.9690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 245.7690 0.0000 245.9690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 245.7690 0.0000 245.9690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 245.7690 0.0000 245.9690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 245.7690 0.0000 245.9690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[50]

  PIN I[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 245.0840 0.0000 245.2840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 245.0840 0.0000 245.2840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 245.0840 0.0000 245.2840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 245.0840 0.0000 245.2840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 245.0840 0.0000 245.2840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[50]

  PIN I[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 246.4520 0.0000 246.6520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 246.4520 0.0000 246.6520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 246.4520 0.0000 246.6520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 246.4520 0.0000 246.6520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 246.4520 0.0000 246.6520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[51]

  PIN O[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 243.0330 0.0000 243.2330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 243.0330 0.0000 243.2330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 243.0330 0.0000 243.2330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 243.0330 0.0000 243.2330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 243.0330 0.0000 243.2330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[48]

  PIN I[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 290.2280 0.0000 290.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 290.2280 0.0000 290.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 290.2280 0.0000 290.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 290.2280 0.0000 290.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 290.2280 0.0000 290.4280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[83]

  PIN O[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 300.4890 0.0000 300.6890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 300.4890 0.0000 300.6890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 300.4890 0.0000 300.6890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 300.4890 0.0000 300.6890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 300.4890 0.0000 300.6890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[90]

  PIN I[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 299.8040 0.0000 300.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 299.8040 0.0000 300.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 299.8040 0.0000 300.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 299.8040 0.0000 300.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 299.8040 0.0000 300.0040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[90]

  PIN I[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 301.1720 0.0000 301.3720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 301.1720 0.0000 301.3720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 301.1720 0.0000 301.3720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 301.1720 0.0000 301.3720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 301.1720 0.0000 301.3720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[91]

  PIN O[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 301.8570 0.0000 302.0570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 301.8570 0.0000 302.0570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 301.8570 0.0000 302.0570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 301.8570 0.0000 302.0570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 301.8570 0.0000 302.0570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[91]

  PIN I[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 295.7000 0.0000 295.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 295.7000 0.0000 295.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 295.7000 0.0000 295.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 295.7000 0.0000 295.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 295.7000 0.0000 295.9000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[87]

  PIN O[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 295.0170 0.0000 295.2170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 295.0170 0.0000 295.2170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 295.0170 0.0000 295.2170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 295.0170 0.0000 295.2170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 295.0170 0.0000 295.2170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[86]

  PIN I[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 297.0680 0.0000 297.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 297.0680 0.0000 297.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 297.0680 0.0000 297.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 297.0680 0.0000 297.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 297.0680 0.0000 297.2680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[88]

  PIN O[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 296.3850 0.0000 296.5850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 296.3850 0.0000 296.5850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 296.3850 0.0000 296.5850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 296.3850 0.0000 296.5850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 296.3850 0.0000 296.5850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[87]

  PIN O[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 297.7530 0.0000 297.9530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 297.7530 0.0000 297.9530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 297.7530 0.0000 297.9530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 297.7530 0.0000 297.9530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 297.7530 0.0000 297.9530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[88]

  PIN O[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 299.1210 0.0000 299.3210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 299.1210 0.0000 299.3210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 299.1210 0.0000 299.3210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 299.1210 0.0000 299.3210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 299.1210 0.0000 299.3210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[89]

  PIN I[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 298.4360 0.0000 298.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 298.4360 0.0000 298.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 298.4360 0.0000 298.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 298.4360 0.0000 298.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 298.4360 0.0000 298.6360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[89]

  PIN I[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 294.3320 0.0000 294.5320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 294.3320 0.0000 294.5320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 294.3320 0.0000 294.5320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 294.3320 0.0000 294.5320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 294.3320 0.0000 294.5320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[86]

  PIN O[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 292.2810 0.0000 292.4810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 292.2810 0.0000 292.4810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 292.2810 0.0000 292.4810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 292.2810 0.0000 292.4810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 292.2810 0.0000 292.4810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[84]

  PIN O[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 290.9130 0.0000 291.1130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 290.9130 0.0000 291.1130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 290.9130 0.0000 291.1130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 290.9130 0.0000 291.1130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 290.9130 0.0000 291.1130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[83]

  PIN I[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 292.9640 0.0000 293.1640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 292.9640 0.0000 293.1640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 292.9640 0.0000 293.1640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 292.9640 0.0000 293.1640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 292.9640 0.0000 293.1640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[85]

  PIN I[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 291.5960 0.0000 291.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 291.5960 0.0000 291.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 291.5960 0.0000 291.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 291.5960 0.0000 291.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 291.5960 0.0000 291.7960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[84]

  PIN O[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 293.6490 0.0000 293.8490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 293.6490 0.0000 293.8490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 293.6490 0.0000 293.8490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 293.6490 0.0000 293.8490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 293.6490 0.0000 293.8490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[85]

  PIN I[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 288.8600 0.0000 289.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 288.8600 0.0000 289.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 288.8600 0.0000 289.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 288.8600 0.0000 289.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 288.8600 0.0000 289.0600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[82]

  PIN O[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 289.5450 0.0000 289.7450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 289.5450 0.0000 289.7450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 289.5450 0.0000 289.7450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 289.5450 0.0000 289.7450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 289.5450 0.0000 289.7450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[82]

  PIN I[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 314.8520 0.0000 315.0520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 314.8520 0.0000 315.0520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 314.8520 0.0000 315.0520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 314.8520 0.0000 315.0520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 314.8520 0.0000 315.0520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[101]

  PIN O[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 311.4330 0.0000 311.6330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 311.4330 0.0000 311.6330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 311.4330 0.0000 311.6330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 311.4330 0.0000 311.6330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 311.4330 0.0000 311.6330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[98]

  PIN I[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 312.1160 0.0000 312.3160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 312.1160 0.0000 312.3160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 312.1160 0.0000 312.3160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 312.1160 0.0000 312.3160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 312.1160 0.0000 312.3160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[99]

  PIN I[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 313.4840 0.0000 313.6840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 313.4840 0.0000 313.6840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 313.4840 0.0000 313.6840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 313.4840 0.0000 313.6840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 313.4840 0.0000 313.6840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[100]

  PIN O[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 312.8010 0.0000 313.0010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 312.8010 0.0000 313.0010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 312.8010 0.0000 313.0010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 312.8010 0.0000 313.0010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 312.8010 0.0000 313.0010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[99]

  PIN O[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 310.0650 0.0000 310.2650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 310.0650 0.0000 310.2650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 310.0650 0.0000 310.2650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 310.0650 0.0000 310.2650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 310.0650 0.0000 310.2650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[97]

  PIN I[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 310.7480 0.0000 310.9480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 310.7480 0.0000 310.9480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 310.7480 0.0000 310.9480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 310.7480 0.0000 310.9480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 310.7480 0.0000 310.9480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[98]

  PIN O[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 308.6970 0.0000 308.8970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 308.6970 0.0000 308.8970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 308.6970 0.0000 308.8970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 308.6970 0.0000 308.8970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 308.6970 0.0000 308.8970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[96]

  PIN I[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 309.3800 0.0000 309.5800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 309.3800 0.0000 309.5800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 309.3800 0.0000 309.5800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 309.3800 0.0000 309.5800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 309.3800 0.0000 309.5800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[97]

  PIN I[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 308.0120 0.0000 308.2120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 308.0120 0.0000 308.2120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 308.0120 0.0000 308.2120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 308.0120 0.0000 308.2120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 308.0120 0.0000 308.2120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[96]

  PIN O[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 307.3290 0.0000 307.5290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 307.3290 0.0000 307.5290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 307.3290 0.0000 307.5290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 307.3290 0.0000 307.5290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 307.3290 0.0000 307.5290 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[95]

  PIN I[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 306.6440 0.0000 306.8440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 306.6440 0.0000 306.8440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 306.6440 0.0000 306.8440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 306.6440 0.0000 306.8440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 306.6440 0.0000 306.8440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[95]

  PIN O[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 305.9610 0.0000 306.1610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 305.9610 0.0000 306.1610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 305.9610 0.0000 306.1610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 305.9610 0.0000 306.1610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 305.9610 0.0000 306.1610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[94]

  PIN I[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 305.2760 0.0000 305.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 305.2760 0.0000 305.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 305.2760 0.0000 305.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 305.2760 0.0000 305.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 305.2760 0.0000 305.4760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[94]

  PIN O[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 304.5930 0.0000 304.7930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 304.5930 0.0000 304.7930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 304.5930 0.0000 304.7930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 304.5930 0.0000 304.7930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 304.5930 0.0000 304.7930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[93]

  PIN O[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 303.2250 0.0000 303.4250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 303.2250 0.0000 303.4250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 303.2250 0.0000 303.4250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 303.2250 0.0000 303.4250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 303.2250 0.0000 303.4250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[92]

  PIN I[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 302.5400 0.0000 302.7400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 302.5400 0.0000 302.7400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 302.5400 0.0000 302.7400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 302.5400 0.0000 302.7400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 302.5400 0.0000 302.7400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[92]

  PIN I[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 303.9080 0.0010 304.1080 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 303.9080 0.0010 304.1080 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 303.9080 0.0000 304.1080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 303.9080 0.0000 304.1080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 303.9080 0.0000 304.1080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[93]

  PIN I[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 328.5320 0.0000 328.7320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 328.5320 0.0000 328.7320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 328.5320 0.0000 328.7320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 328.5320 0.0000 328.7320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 328.5320 0.0000 328.7320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[111]

  PIN O[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 326.4810 0.0000 326.6810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 326.4810 0.0000 326.6810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 326.4810 0.0000 326.6810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 326.4810 0.0000 326.6810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 326.4810 0.0000 326.6810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[109]

  PIN I[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 325.7960 0.0000 325.9960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 325.7960 0.0000 325.9960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 325.7960 0.0000 325.9960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 325.7960 0.0000 325.9960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 325.7960 0.0000 325.9960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[109]

  PIN O[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 323.7450 0.0000 323.9450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 323.7450 0.0000 323.9450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 323.7450 0.0000 323.9450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 323.7450 0.0000 323.9450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 323.7450 0.0000 323.9450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[107]

  PIN I[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 324.4280 0.0000 324.6280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 324.4280 0.0000 324.6280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 324.4280 0.0000 324.6280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 324.4280 0.0000 324.6280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 324.4280 0.0000 324.6280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[108]

  PIN O[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 325.1130 0.0000 325.3130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 325.1130 0.0000 325.3130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 325.1130 0.0000 325.3130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 325.1130 0.0000 325.3130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 325.1130 0.0000 325.3130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[108]

  PIN I[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 321.6920 0.0000 321.8920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 321.6920 0.0000 321.8920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 321.6920 0.0000 321.8920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 321.6920 0.0000 321.8920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 321.6920 0.0000 321.8920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[106]

  PIN I[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 323.0600 0.0000 323.2600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 323.0600 0.0000 323.2600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 323.0600 0.0000 323.2600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 323.0600 0.0000 323.2600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 323.0600 0.0000 323.2600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[107]

  PIN O[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 322.3770 0.0000 322.5770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 322.3770 0.0000 322.5770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 322.3770 0.0000 322.5770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 322.3770 0.0000 322.5770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 322.3770 0.0000 322.5770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[106]

  PIN O[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 321.0090 0.0000 321.2090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 321.0090 0.0000 321.2090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 321.0090 0.0000 321.2090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 321.0090 0.0000 321.2090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 321.0090 0.0000 321.2090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[105]

  PIN O[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 319.6410 0.0000 319.8410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 319.6410 0.0000 319.8410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 319.6410 0.0000 319.8410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 319.6410 0.0000 319.8410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 319.6410 0.0000 319.8410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[104]

  PIN I[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 318.9560 0.0000 319.1560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 318.9560 0.0000 319.1560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 318.9560 0.0000 319.1560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 318.9560 0.0000 319.1560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 318.9560 0.0000 319.1560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[104]

  PIN I[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 320.3240 0.0000 320.5240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 320.3240 0.0000 320.5240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 320.3240 0.0000 320.5240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 320.3240 0.0000 320.5240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 320.3240 0.0000 320.5240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[105]

  PIN O[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 318.2730 0.0000 318.4730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 318.2730 0.0000 318.4730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 318.2730 0.0000 318.4730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 318.2730 0.0000 318.4730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 318.2730 0.0000 318.4730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[103]

  PIN I[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 317.5880 0.0000 317.7880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 317.5880 0.0000 317.7880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 317.5880 0.0000 317.7880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 317.5880 0.0000 317.7880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 317.5880 0.0000 317.7880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[103]

  PIN O[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 316.9050 0.0000 317.1050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 316.9050 0.0000 317.1050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 316.9050 0.0000 317.1050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 316.9050 0.0000 317.1050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 316.9050 0.0000 317.1050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[102]

  PIN I[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 316.2200 0.0000 316.4200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 316.2200 0.0000 316.4200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 316.2200 0.0000 316.4200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 316.2200 0.0000 316.4200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 316.2200 0.0000 316.4200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[102]

  PIN O[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 314.1690 0.0000 314.3690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 314.1690 0.0000 314.3690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 314.1690 0.0000 314.3690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 314.1690 0.0000 314.3690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 314.1690 0.0000 314.3690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[100]

  PIN O[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 315.5370 0.0000 315.7370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 315.5370 0.0000 315.7370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 315.5370 0.0000 315.7370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 315.5370 0.0000 315.7370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 315.5370 0.0000 315.7370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[101]

  PIN I[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 340.8440 0.0000 341.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 340.8440 0.0000 341.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 340.8440 0.0000 341.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 340.8440 0.0000 341.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 340.8440 0.0000 341.0440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[120]

  PIN I[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 339.4760 0.0000 339.6760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 339.4760 0.0000 339.6760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 339.4760 0.0000 339.6760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 339.4760 0.0000 339.6760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 339.4760 0.0000 339.6760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[119]

  PIN O[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 340.1610 0.0000 340.3610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 340.1610 0.0000 340.3610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 340.1610 0.0000 340.3610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 340.1610 0.0000 340.3610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 340.1610 0.0000 340.3610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[119]

  PIN I[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 336.7400 0.0000 336.9400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 336.7400 0.0000 336.9400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 336.7400 0.0000 336.9400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 336.7400 0.0000 336.9400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 336.7400 0.0000 336.9400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[117]

  PIN O[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 337.4250 0.0000 337.6250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 337.4250 0.0000 337.6250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 337.4250 0.0000 337.6250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 337.4250 0.0000 337.6250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 337.4250 0.0000 337.6250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[117]

  PIN I[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 334.0040 0.0000 334.2040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 334.0040 0.0000 334.2040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 334.0040 0.0000 334.2040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 334.0040 0.0000 334.2040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 334.0040 0.0000 334.2040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[115]

  PIN O[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 334.6890 0.0000 334.8890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 334.6890 0.0000 334.8890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 334.6890 0.0000 334.8890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 334.6890 0.0000 334.8890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 334.6890 0.0000 334.8890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[115]

  PIN I[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 335.3720 0.0000 335.5720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 335.3720 0.0000 335.5720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 335.3720 0.0000 335.5720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 335.3720 0.0000 335.5720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 335.3720 0.0000 335.5720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[116]

  PIN O[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 336.0570 0.0000 336.2570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 336.0570 0.0000 336.2570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 336.0570 0.0000 336.2570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 336.0570 0.0000 336.2570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 336.0570 0.0000 336.2570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[116]

  PIN I[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 331.2680 0.0000 331.4680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 331.2680 0.0000 331.4680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 331.2680 0.0000 331.4680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 331.2680 0.0000 331.4680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 331.2680 0.0000 331.4680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[113]

  PIN O[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 330.5850 0.0000 330.7850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 330.5850 0.0000 330.7850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 330.5850 0.0000 330.7850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 330.5850 0.0000 330.7850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 330.5850 0.0000 330.7850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[112]

  PIN I[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 332.6360 0.0000 332.8360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 332.6360 0.0000 332.8360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 332.6360 0.0000 332.8360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 332.6360 0.0000 332.8360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 332.6360 0.0000 332.8360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[114]

  PIN I[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 329.9000 0.0000 330.1000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 329.9000 0.0000 330.1000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 329.9000 0.0000 330.1000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 329.9000 0.0000 330.1000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 329.9000 0.0000 330.1000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[112]

  PIN O[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 331.9530 0.0000 332.1530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 331.9530 0.0000 332.1530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 331.9530 0.0000 332.1530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 331.9530 0.0000 332.1530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 331.9530 0.0000 332.1530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[113]

  PIN O[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 333.3210 0.0000 333.5210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 333.3210 0.0000 333.5210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 333.3210 0.0000 333.5210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 333.3210 0.0000 333.5210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 333.3210 0.0000 333.5210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[114]

  PIN O[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 327.8490 0.0000 328.0490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 327.8490 0.0000 328.0490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 327.8490 0.0000 328.0490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 327.8490 0.0000 328.0490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 327.8490 0.0000 328.0490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[110]

  PIN I[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 327.1640 0.0000 327.3640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 327.1640 0.0000 327.3640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 327.1640 0.0000 327.3640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 327.1640 0.0000 327.3640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 327.1640 0.0000 327.3640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[110]

  PIN O[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 329.2170 0.0000 329.4170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 329.2170 0.0000 329.4170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 329.2170 0.0000 329.4170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 329.2170 0.0000 329.4170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 329.2170 0.0000 329.4170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[111]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 17.2900 372.8790 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 17.2900 372.8790 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 17.2900 372.8790 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 17.2900 372.8790 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 17.2900 372.8790 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 372.6790 16.8280 372.8790 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 372.6790 16.8280 372.8790 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 372.6790 16.8280 372.8790 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 372.6790 16.8280 372.8790 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 372.6790 16.8280 372.8790 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN O[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 349.7370 0.0000 349.9370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 349.7370 0.0000 349.9370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 349.7370 0.0000 349.9370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 349.7370 0.0000 349.9370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 349.7370 0.0000 349.9370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[126]
  OBS
    LAYER M2 ;
      RECT 0.0000 292.3480 372.8790 309.2530 ;
      RECT 0.0000 272.9310 371.9850 309.2530 ;
      RECT 0.0000 0.0000 175.9840 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 287.1530 371.9850 292.3480 ;
      RECT 0.0000 272.9310 372.8790 287.1530 ;
      RECT 0.0000 271.3310 371.9790 272.9310 ;
      RECT 371.3780 289.0960 372.8790 290.7480 ;
      RECT 0.0000 265.7010 372.8790 271.3310 ;
      RECT 0.0000 262.5110 371.9790 265.7010 ;
      RECT 0.0000 256.8810 372.8790 262.5110 ;
      RECT 0.0000 253.6910 371.9790 256.8810 ;
      RECT 0.0000 248.0650 372.8790 253.6910 ;
      RECT 0.0000 244.8750 371.9790 248.0650 ;
      RECT 0.0000 95.0160 372.8790 244.8750 ;
      RECT 0.0000 93.4160 371.9790 95.0160 ;
      RECT 0.0000 18.1900 372.8790 93.4160 ;
      RECT 0.0000 16.1280 371.9790 18.1900 ;
      RECT 0.0000 10.7200 372.8790 16.1280 ;
      RECT 0.0000 9.1200 371.9790 10.7200 ;
      RECT 0.0000 0.9000 372.8790 9.1200 ;
      RECT 0.0000 0.0000 175.9840 0.9000 ;
      RECT 352.6780 0.0000 372.8790 9.1200 ;
      RECT 352.6780 0.0000 372.8790 0.9000 ;
    LAYER M1 ;
      RECT 372.0790 246.3750 372.8790 246.5650 ;
      RECT 372.0790 255.1910 372.8790 255.3810 ;
      RECT 372.0790 264.0110 372.8790 264.2010 ;
      RECT 371.3780 288.9960 372.8790 290.8480 ;
      RECT 0.0000 265.6010 372.8790 271.4310 ;
      RECT 0.0000 262.6110 372.0790 265.6010 ;
      RECT 0.0000 256.7810 372.8790 262.6110 ;
      RECT 0.0000 253.7910 372.0790 256.7810 ;
      RECT 0.0000 247.9650 372.8790 253.7910 ;
      RECT 0.0000 244.9750 372.0790 247.9650 ;
      RECT 0.0000 94.9160 372.8790 244.9750 ;
      RECT 0.0000 93.5160 372.0790 94.9160 ;
      RECT 0.0000 18.0900 372.8790 93.5160 ;
      RECT 0.0000 16.2280 372.0790 18.0900 ;
      RECT 0.0000 10.6200 372.8790 16.2280 ;
      RECT 0.0000 9.2200 372.0790 10.6200 ;
      RECT 0.0000 0.8000 372.8790 9.2200 ;
      RECT 0.0000 0.0000 176.0840 0.8000 ;
      RECT 352.5780 0.0000 372.8790 9.2200 ;
      RECT 352.5780 0.0000 372.8790 0.8000 ;
      RECT 0.0000 292.2480 372.8790 309.2530 ;
      RECT 0.0000 272.8310 372.0850 309.2530 ;
      RECT 0.0000 0.0000 176.0840 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 0.8000 372.0790 309.2530 ;
      RECT 0.0000 287.2530 372.0850 292.2480 ;
      RECT 0.0000 272.8310 372.8790 287.2530 ;
      RECT 0.0000 271.4310 372.0790 272.8310 ;
    LAYER PO ;
      RECT 0.0000 0.0000 372.8790 309.2530 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 372.8790 309.2530 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 372.8790 309.2530 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 372.8790 309.2530 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 372.8790 309.2530 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 372.8790 309.2530 ;
    LAYER M5 ;
      RECT 372.2890 308.2530 372.8790 309.2530 ;
      RECT 371.3780 289.0960 372.8790 290.7480 ;
      RECT 0.0000 0.0000 175.9840 0.9000 ;
      RECT 352.6780 0.0000 372.8790 0.9000 ;
      RECT 0.0000 265.7010 372.8790 271.3310 ;
      RECT 0.0000 262.5110 371.9790 265.7010 ;
      RECT 0.0000 256.8810 372.8790 262.5110 ;
      RECT 0.0000 253.6910 371.9790 256.8810 ;
      RECT 0.0000 248.0650 372.8790 253.6910 ;
      RECT 0.0000 244.8750 371.9790 248.0650 ;
      RECT 0.0000 95.0160 372.8790 244.8750 ;
      RECT 0.0000 93.4160 371.9790 95.0160 ;
      RECT 0.0000 18.1900 372.8790 93.4160 ;
      RECT 0.0000 16.1280 371.9790 18.1900 ;
      RECT 0.0000 10.7200 372.8790 16.1280 ;
      RECT 0.0000 9.1200 371.9790 10.7200 ;
      RECT 0.0000 0.9010 372.8790 9.1200 ;
      RECT 0.0000 0.9000 177.3520 0.9010 ;
      RECT 178.9520 0.9000 240.2800 0.9010 ;
      RECT 241.8800 0.9000 303.2080 0.9010 ;
      RECT 304.8080 0.9000 372.8790 9.1200 ;
      RECT 304.8080 0.9000 372.8790 0.9010 ;
      RECT 352.6780 0.0000 372.8790 9.1200 ;
      RECT 0.0000 0.9000 177.3520 308.2530 ;
      RECT 0.0000 292.3480 372.8790 308.2530 ;
      RECT 0.0000 272.9310 371.9850 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 0.9010 371.9790 308.2530 ;
      RECT 0.0000 287.1530 371.9850 292.3480 ;
      RECT 0.0000 272.9310 372.8790 287.1530 ;
      RECT 0.0000 271.3310 371.9790 272.9310 ;
      RECT 178.9520 0.9000 240.2800 308.2530 ;
      RECT 241.8800 0.9000 303.2080 308.2530 ;
    LAYER M4 ;
      RECT 371.3780 289.0960 372.8790 290.7480 ;
      RECT 0.0000 0.0000 175.9840 0.9000 ;
      RECT 352.6780 0.0000 372.8790 0.9000 ;
      RECT 0.0000 265.7010 372.8790 271.3310 ;
      RECT 0.0000 262.5110 371.9790 265.7010 ;
      RECT 0.0000 256.8810 372.8790 262.5110 ;
      RECT 0.0000 253.6910 371.9790 256.8810 ;
      RECT 0.0000 248.0650 372.8790 253.6910 ;
      RECT 0.0000 244.8750 371.9790 248.0650 ;
      RECT 0.0000 95.0160 372.8790 244.8750 ;
      RECT 0.0000 93.4160 371.9790 95.0160 ;
      RECT 0.0000 18.1900 372.8790 93.4160 ;
      RECT 0.0000 16.1280 371.9790 18.1900 ;
      RECT 0.0000 10.7200 372.8790 16.1280 ;
      RECT 0.0000 9.1200 371.9790 10.7200 ;
      RECT 0.0000 0.9010 372.8790 9.1200 ;
      RECT 0.0000 0.9000 177.3520 0.9010 ;
      RECT 178.9520 0.9000 240.2800 0.9010 ;
      RECT 241.8800 0.9000 303.2080 0.9010 ;
      RECT 304.8080 0.9000 372.8790 9.1200 ;
      RECT 304.8080 0.9000 372.8790 0.9010 ;
      RECT 352.6780 0.0000 372.8790 9.1200 ;
      RECT 0.0000 0.9000 177.3520 309.2530 ;
      RECT 0.0000 292.3480 372.8790 309.2530 ;
      RECT 0.0000 272.9310 371.9850 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 0.9010 371.9790 309.2530 ;
      RECT 0.0000 287.1530 371.9850 292.3480 ;
      RECT 0.0000 272.9310 372.8790 287.1530 ;
      RECT 0.0000 271.3310 371.9790 272.9310 ;
      RECT 178.9520 0.9000 240.2800 309.2530 ;
      RECT 241.8800 0.9000 303.2080 309.2530 ;
    LAYER M3 ;
      RECT 371.3780 289.0960 372.8790 290.7480 ;
      RECT 0.0000 265.7010 372.8790 271.3310 ;
      RECT 0.0000 262.5110 371.9790 265.7010 ;
      RECT 0.0000 256.8810 372.8790 262.5110 ;
      RECT 0.0000 253.6910 371.9790 256.8810 ;
      RECT 0.0000 248.0650 372.8790 253.6910 ;
      RECT 0.0000 244.8750 371.9790 248.0650 ;
      RECT 0.0000 95.0160 372.8790 244.8750 ;
      RECT 0.0000 93.4160 371.9790 95.0160 ;
      RECT 0.0000 18.1900 372.8790 93.4160 ;
      RECT 0.0000 16.1280 371.9790 18.1900 ;
      RECT 0.0000 10.7200 372.8790 16.1280 ;
      RECT 0.0000 9.1200 371.9790 10.7200 ;
      RECT 0.0000 0.9000 372.8790 9.1200 ;
      RECT 0.0000 0.0000 175.9840 0.9000 ;
      RECT 352.6780 0.0000 372.8790 9.1200 ;
      RECT 352.6780 0.0000 372.8790 0.9000 ;
      RECT 0.0000 292.3480 372.8790 309.2530 ;
      RECT 0.0000 272.9310 371.9850 309.2530 ;
      RECT 0.0000 0.0000 175.9840 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 0.9000 371.9790 309.2530 ;
      RECT 0.0000 287.1530 371.9850 292.3480 ;
      RECT 0.0000 272.9310 372.8790 287.1530 ;
      RECT 0.0000 271.3310 371.9790 272.9310 ;
  END
END SRAMLP1RW256x128

MACRO SRAMLP1RW512x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 59.822 BY 244.564 ;
  SYMMETRY X Y R90 ;

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6250 182.3150 59.8220 182.5150 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6250 182.3150 59.8220 182.5150 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6250 182.3150 59.8220 182.5150 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6250 182.3150 59.8220 182.5150 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6250 182.3150 59.8220 182.5150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.305828 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.305828 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16906 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16906 LAYER M2 ;
    ANTENNAMAXAREACAR 12.97459 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[5]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.5170 0.0000 34.7170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.5170 0.0000 34.7170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.5170 0.0000 34.7170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.5170 0.0000 34.7170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.5170 0.0000 34.7170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.917257 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.917257 LAYER M2 ;
    ANTENNAMAXAREACAR 7.362508 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.52312 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52312 LAYER M3 ;
    ANTENNAMAXAREACAR 11.01034 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 17.9100 59.8220 18.1100 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 17.9100 59.8220 18.1100 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 17.9100 59.8220 18.1100 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 17.9100 59.8220 18.1100 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 17.9100 59.8220 18.1100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.49402 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.49402 LAYER M2 ;
    ANTENNAGATEAREA 21.3756 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 518.989 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 518.989 LAYER M3 ;
    ANTENNAMAXAREACAR 10779.46 LAYER M3 ;
    ANTENNAGATEAREA 21.3756 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 2003.716 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2003.716 LAYER M4 ;
    ANTENNAMAXAREACAR 10873.2 LAYER M4 ;
    ANTENNAGATEAREA 21.3756 LAYER M5 ;
    ANTENNAGATEAREA 21.3756 LAYER M6 ;
    ANTENNAGATEAREA 21.3756 LAYER M7 ;
    ANTENNAGATEAREA 21.3756 LAYER M8 ;
    ANTENNAGATEAREA 21.3756 LAYER M9 ;
    ANTENNAGATEAREA 21.3756 LAYER MRDL ;
  END CSB

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 9.7780 59.8220 9.9780 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 9.7780 59.8220 9.9780 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 9.7780 59.8220 9.9780 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 9.7780 59.8220 9.9780 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 9.7780 59.8220 9.9780 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.839697 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.839697 LAYER M2 ;
    ANTENNAMAXAREACAR 13.63038 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.52312 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52312 LAYER M3 ;
    ANTENNAMAXAREACAR 17.21068 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.52312 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52312 LAYER M4 ;
    ANTENNAMAXAREACAR 20.79091 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 21.82718 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 48.1710 244.2630 48.4710 244.5630 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.0700 244.2630 49.3700 244.5630 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.9710 244.2630 50.2710 244.5630 ;
    END
  END VDDL

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 29.4170 59.8220 29.6170 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 29.4170 59.8220 29.6170 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 29.4170 59.8220 29.6170 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 29.4170 59.8220 29.6170 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 29.4170 59.8220 29.6170 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.32691 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.32691 LAYER M2 ;
  END A[7]

  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 28.6920 59.8220 28.8920 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 28.6920 59.8220 28.8920 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 28.6920 59.8220 28.8920 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 28.6920 59.8220 28.8920 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 28.6920 59.8220 28.8920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M2 ;
  END A[8]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5800 0.0000 23.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5800 0.0000 23.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5800 0.0000 23.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5800 0.0000 23.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5800 0.0000 23.7800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 1.5102 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 24.81794 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.81794 LAYER M3 ;
    ANTENNAMAXAREACAR 57.43748 LAYER M3 ;
    ANTENNAGATEAREA 3.4446 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 76.69425 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 76.69425 LAYER M4 ;
    ANTENNAMAXAREACAR 36.63142 LAYER M4 ;
    ANTENNAGATEAREA 31.9764 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 9514.22 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 9514.22 LAYER M5 ;
    ANTENNAMAXAREACAR 328.049 LAYER M5 ;
    ANTENNAGATEAREA 31.9764 LAYER M6 ;
    ANTENNAGATEAREA 31.9764 LAYER M7 ;
    ANTENNAGATEAREA 31.9764 LAYER M8 ;
    ANTENNAGATEAREA 31.9764 LAYER M9 ;
    ANTENNAGATEAREA 31.9764 LAYER MRDL ;
  END I[0]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6140 0.0000 25.8140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6140 0.0000 25.8140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6140 0.0000 25.8140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6140 0.0000 25.8140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6140 0.0000 25.8140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[7]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6230 191.1330 59.8220 191.3330 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6230 191.1330 59.8220 191.3330 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6230 191.1330 59.8220 191.3330 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6230 191.1330 59.8220 191.3330 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6230 191.1330 59.8220 191.3330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.306008 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.306008 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16934 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16934 LAYER M2 ;
    ANTENNAMAXAREACAR 12.98716 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[3]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 180.7490 59.8220 180.9490 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 180.7490 59.8220 180.9490 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 180.7490 59.8220 180.9490 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 180.7490 59.8220 180.9490 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 180.7490 59.8220 180.9490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.306198 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.306198 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M2 ;
    ANTENNAMAXAREACAR 12.99617 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[6]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7880 0.0000 31.9880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7880 0.0000 31.9880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7880 0.0000 31.9880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7880 0.0000 31.9880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7880 0.0000 31.9880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[3]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1560 0.0000 33.3560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1560 0.0000 33.3560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1560 0.0000 33.3560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1560 0.0000 33.3560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1560 0.0000 33.3560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[5]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2460 0.0000 24.4460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2460 0.0000 24.4460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2460 0.0000 24.4460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2460 0.0000 24.4460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2460 0.0000 24.4460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[0]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0910 0.0000 31.2910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0910 0.0000 31.2910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0910 0.0000 31.2910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0910 0.0000 31.2910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0910 0.0000 31.2910 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[2]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4510 0.0000 32.6510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4510 0.0000 32.6510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4510 0.0000 32.6510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4510 0.0000 32.6510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4510 0.0000 32.6510 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[3]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.3160 0.0000 26.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.3160 0.0000 26.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.3160 0.0000 26.5160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.3160 0.0000 26.5160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.3160 0.0000 26.5160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[1]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7170 0.0000 29.9170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7170 0.0000 29.9170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7170 0.0000 29.9170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7170 0.0000 29.9170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7170 0.0000 29.9170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[4]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.9480 0.0000 25.1480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.9480 0.0000 25.1480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.9480 0.0000 25.1480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.9480 0.0000 25.1480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.9480 0.0000 25.1480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[7]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9830 0.0000 27.1830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9830 0.0000 27.1830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9830 0.0000 27.1830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9830 0.0000 27.1830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9830 0.0000 27.1830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[1]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.0520 0.0000 29.2520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.0520 0.0000 29.2520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.0520 0.0000 29.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.0520 0.0000 29.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.0520 0.0000 29.2520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[4]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8080 0.0000 34.0080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8080 0.0000 34.0080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8080 0.0000 34.0080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8080 0.0000 34.0080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8080 0.0000 34.0080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.570708 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.570708 LAYER M3 ;
  END O[5]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 18.6650 59.8220 18.8650 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 18.6650 59.8220 18.8650 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 18.6650 59.8220 18.8650 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 18.6650 59.8220 18.8650 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 18.6650 59.8220 18.8650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.74759 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74759 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M2 ;
    ANTENNAMAXAREACAR 25.05535 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CE

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.4200 0.0000 30.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.4200 0.0000 30.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.4200 0.0000 30.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.4200 0.0000 30.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.4200 0.0000 30.6200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[2]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3530 0.0000 28.5530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3530 0.0000 28.5530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3540 0.0000 28.5540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3540 0.0000 28.5540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3540 0.0000 28.5540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END O[6]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6840 0.0000 27.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6840 0.0000 27.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6840 0.0000 27.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6840 0.0000 27.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6840 0.0000 27.8840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
  END I[6]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6250 189.5700 59.8220 189.7700 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6250 189.5700 59.8220 189.7700 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6250 189.5700 59.8220 189.7700 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6250 189.5700 59.8220 189.7700 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6250 189.5700 59.8220 189.7700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.305828 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.305828 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16906 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16906 LAYER M2 ;
    ANTENNAMAXAREACAR 12.97459 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[4]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6280 227.5670 59.8220 227.7670 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6280 227.5670 59.8220 227.7670 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6280 227.5670 59.8220 227.7670 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6280 227.5670 59.8220 227.7670 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6280 227.5670 59.8220 227.7670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.222445 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.222445 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END LS

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6280 224.4140 59.8220 224.6140 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6280 224.4140 59.8220 224.6140 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6280 224.4140 59.8220 224.6140 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6280 224.4140 59.8220 224.6140 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6280 224.4140 59.8220 224.6140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0213 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.323462 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.323462 LAYER M1 ;
    ANTENNAGATEAREA 2.4783 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 66.29205 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.29205 LAYER M2 ;
    ANTENNAMAXAREACAR 35.42044 LAYER M2 ;
    ANTENNAGATEAREA 2.4783 LAYER M3 ;
    ANTENNAGATEAREA 2.4783 LAYER M4 ;
    ANTENNAGATEAREA 2.4783 LAYER M5 ;
    ANTENNAGATEAREA 2.4783 LAYER M6 ;
    ANTENNAGATEAREA 2.4783 LAYER M7 ;
    ANTENNAGATEAREA 2.4783 LAYER M8 ;
    ANTENNAGATEAREA 2.4783 LAYER M9 ;
    ANTENNAGATEAREA 2.4783 LAYER MRDL ;
  END DS

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6280 223.8530 59.8220 224.0530 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6280 223.8530 59.8220 224.0530 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6280 223.8530 59.8220 224.0530 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6280 223.8530 59.8220 224.0530 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6280 223.8530 59.8220 224.0530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M2 ;
  END SD

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 57.1730 244.2630 57.4720 244.5630 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.0730 244.2630 58.3730 244.5630 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.2720 244.2630 56.5720 244.5630 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 43.2190 244.2640 43.5200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.4180 244.2640 50.7180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.3180 244.2640 51.6180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.2180 244.2640 52.5180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.0180 244.2640 54.3180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.9180 244.2640 55.2180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.8220 244.2640 56.1220 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.6180 244.2640 48.9180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.7180 244.2640 48.0180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.8180 244.2640 47.1180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.0180 244.2640 45.3180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.2190 244.2640 25.5190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.4190 244.2640 23.7190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.5200 244.2640 22.8200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.6200 244.2640 21.9200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.8200 244.2640 20.1200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.9200 244.2640 19.2200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0200 244.2640 18.3200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.2200 244.2640 16.5200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.3200 244.2640 15.6200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.4200 244.2640 14.7200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6200 244.2640 12.9200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.7180 244.2640 57.0180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.1190 244.2640 53.4190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.5190 244.2640 49.8190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.9190 244.2640 46.2190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.1180 244.2640 44.4180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.3200 244.2640 24.6200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.7210 244.2640 21.0210 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1210 244.2640 17.4210 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.5210 244.2640 13.8210 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7200 244.2640 12.0200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.3180 244.2640 42.6170 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.9200 244.2640 10.2190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.9190 244.2640 37.2190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.5210 244.2640 4.8210 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.4190 244.2640 41.7190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.0210 244.2640 9.3210 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.5180 244.2640 40.8180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.1200 244.2640 8.4200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.0180 244.2640 36.3180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6200 244.2640 3.9200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.8180 244.2640 38.1170 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.4200 244.2640 5.7190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.1180 244.2640 35.4180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7200 244.2640 3.0200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.6180 244.2640 39.9180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.2200 244.2640 7.5200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.0190 244.2640 27.3180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.1190 244.2640 26.4190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.2190 244.2640 34.5200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.8210 244.2640 2.1220 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.8180 244.2640 29.1190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.7180 244.2640 30.0190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.9190 244.2640 28.2180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.5180 244.2640 31.8180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.3180 244.2640 33.6170 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.9200 244.2640 1.2190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.4190 244.2640 32.7190 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0210 244.2640 0.3210 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.6180 244.2640 30.9180 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.7190 244.2640 39.0200 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.3210 244.2640 6.6220 244.5640 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.8210 244.2640 11.1220 244.5640 ;
    END
  END VSS

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6250 199.9640 59.8220 200.1640 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6250 199.9640 59.8220 200.1640 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6250 199.9640 59.8220 200.1640 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6250 199.9640 59.8220 200.1640 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6250 199.9640 59.8220 200.1640 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.307353 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.307353 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16906 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16906 LAYER M2 ;
    ANTENNAMAXAREACAR 13.01625 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[1]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6220 207.2540 59.8220 207.4540 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6220 207.2540 59.8220 207.4540 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6220 207.2540 59.8220 207.4540 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6220 207.2540 59.8220 207.4540 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6220 207.2540 59.8220 207.4540 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.306098 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.306098 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16948 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16948 LAYER M2 ;
    ANTENNAMAXAREACAR 12.99344 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[0]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.6380 198.4320 59.8220 198.6320 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.6380 198.4320 59.8220 198.6320 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.6380 198.4320 59.8220 198.6320 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.6380 198.4320 59.8220 198.6320 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.6380 198.4320 59.8220 198.6320 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.307403 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.307403 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.16724 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16724 LAYER M2 ;
    ANTENNAMAXAREACAR 12.96789 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[2]
  OBS
    LAYER M2 ;
      RECT 0.0000 188.8700 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 183.2150 59.8220 188.8700 ;
      RECT 0.0000 181.6490 58.9250 183.2150 ;
      RECT 0.0000 180.0490 58.9220 181.6490 ;
      RECT 0.0000 30.3170 59.8220 180.0490 ;
      RECT 0.0000 27.9920 58.9220 30.3170 ;
      RECT 0.0000 19.5650 59.8220 27.9920 ;
      RECT 0.0000 17.2100 58.9220 19.5650 ;
      RECT 0.0000 10.6780 59.8220 17.2100 ;
      RECT 0.0000 9.0780 58.9220 10.6780 ;
      RECT 0.0000 0.9000 59.8220 9.0780 ;
      RECT 0.0000 0.0000 22.8800 0.9000 ;
      RECT 35.4170 0.0000 59.8220 9.0780 ;
      RECT 35.4170 0.0000 59.8220 0.9000 ;
      RECT 0.0000 228.4670 59.8220 244.5640 ;
      RECT 0.0000 208.1540 58.9280 244.5640 ;
      RECT 0.0000 0.0000 22.8800 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 223.1530 58.9280 228.4670 ;
      RECT 0.0000 208.1540 59.8220 223.1530 ;
      RECT 0.0000 206.5540 58.9220 208.1540 ;
      RECT 58.3210 225.3140 59.8220 226.8670 ;
      RECT 0.0000 200.8640 59.8220 206.5540 ;
      RECT 0.0000 192.0330 58.9250 206.5540 ;
      RECT 0.0000 181.6490 58.9230 206.5540 ;
      RECT 0.0000 199.2640 58.9250 200.8640 ;
      RECT 0.0000 197.7320 58.9380 199.2640 ;
      RECT 0.0000 192.0330 58.9380 199.2640 ;
      RECT 0.0000 192.0330 59.8220 197.7320 ;
      RECT 0.0000 190.4330 58.9230 192.0330 ;
    LAYER M1 ;
      RECT 59.0380 199.2320 59.8220 199.3640 ;
      RECT 59.0250 181.5490 59.8220 181.7150 ;
      RECT 59.0250 190.3700 59.8220 190.5330 ;
      RECT 58.3210 225.2140 59.8220 226.9670 ;
      RECT 0.0000 200.7640 59.8220 206.6540 ;
      RECT 0.0000 191.9330 59.0250 206.6540 ;
      RECT 0.0000 181.5490 59.0230 206.6540 ;
      RECT 0.0000 199.3640 59.0250 200.7640 ;
      RECT 0.0000 197.8320 59.0380 199.3640 ;
      RECT 0.0000 191.9330 59.0380 199.3640 ;
      RECT 0.0000 191.9330 59.8220 197.8320 ;
      RECT 0.0000 190.5330 59.0230 191.9330 ;
      RECT 0.0000 188.9700 59.0250 190.5330 ;
      RECT 0.0000 181.5490 59.0250 190.5330 ;
      RECT 0.0000 181.5490 59.0250 190.5330 ;
      RECT 0.0000 183.1150 59.8220 188.9700 ;
      RECT 0.0000 181.5490 59.0250 183.1150 ;
      RECT 0.0000 180.1490 59.0220 181.5490 ;
      RECT 0.0000 30.2170 59.8220 180.1490 ;
      RECT 0.0000 28.0920 59.0220 30.2170 ;
      RECT 0.0000 19.4650 59.8220 28.0920 ;
      RECT 0.0000 17.3100 59.0220 19.4650 ;
      RECT 0.0000 10.5780 59.8220 17.3100 ;
      RECT 0.0000 9.1780 59.0220 10.5780 ;
      RECT 0.0000 0.8000 59.8220 9.1780 ;
      RECT 0.0000 0.0000 22.9800 0.8000 ;
      RECT 35.3170 0.0000 59.8220 9.1780 ;
      RECT 35.3170 0.0000 59.8220 0.8000 ;
      RECT 0.0000 228.3670 59.8220 244.5640 ;
      RECT 0.0000 208.0540 59.0280 244.5640 ;
      RECT 0.0000 0.0000 22.9800 244.5640 ;
      RECT 0.0000 0.8000 59.0220 244.5640 ;
      RECT 0.0000 0.8000 59.0220 244.5640 ;
      RECT 0.0000 0.8000 59.0220 244.5640 ;
      RECT 0.0000 0.8000 59.0220 244.5640 ;
      RECT 0.0000 0.8000 59.0220 244.5640 ;
      RECT 0.0000 223.2530 59.0280 228.3670 ;
      RECT 0.0000 208.0540 59.8220 223.2530 ;
      RECT 0.0000 206.6540 59.0220 208.0540 ;
    LAYER PO ;
      RECT 0.0000 0.0000 59.8220 244.5640 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 59.8220 244.5640 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 59.8220 244.5640 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 59.8220 244.5640 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 59.8220 244.5640 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 59.8220 244.5640 ;
    LAYER M5 ;
      RECT 59.0730 243.5630 59.8220 244.5640 ;
      RECT 58.3210 225.3140 59.8220 226.8670 ;
      RECT 50.9710 243.5630 55.5720 243.5640 ;
      RECT 50.9710 0.9000 55.5720 243.5640 ;
      RECT 0.0000 243.5630 47.4710 243.5640 ;
      RECT 0.0000 0.9000 47.4710 243.5640 ;
      RECT 0.0000 0.0000 22.8800 243.5630 ;
      RECT 0.0000 228.4670 59.8220 243.5630 ;
      RECT 0.0000 208.1540 58.9280 243.5630 ;
      RECT 0.0000 0.9000 58.9220 243.5630 ;
      RECT 0.0000 0.9000 58.9220 243.5630 ;
      RECT 0.0000 0.9000 58.9220 243.5630 ;
      RECT 0.0000 0.9000 58.9220 243.5630 ;
      RECT 0.0000 0.9000 58.9220 243.5630 ;
      RECT 0.0000 223.1530 58.9280 228.4670 ;
      RECT 0.0000 208.1540 59.8220 223.1530 ;
      RECT 0.0000 206.5540 58.9220 208.1540 ;
      RECT 0.0000 200.8640 59.8220 206.5540 ;
      RECT 0.0000 192.0330 58.9250 206.5540 ;
      RECT 0.0000 181.6490 58.9230 206.5540 ;
      RECT 0.0000 199.2640 58.9250 200.8640 ;
      RECT 0.0000 197.7320 58.9380 199.2640 ;
      RECT 0.0000 192.0330 58.9380 199.2640 ;
      RECT 0.0000 192.0330 59.8220 197.7320 ;
      RECT 0.0000 190.4330 58.9230 192.0330 ;
      RECT 0.0000 188.8700 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 183.2150 59.8220 188.8700 ;
      RECT 0.0000 181.6490 58.9250 183.2150 ;
      RECT 0.0000 180.0490 58.9220 181.6490 ;
      RECT 0.0000 30.3170 59.8220 180.0490 ;
      RECT 0.0000 27.9920 58.9220 30.3170 ;
      RECT 0.0000 19.5650 59.8220 27.9920 ;
      RECT 0.0000 17.2100 58.9220 19.5650 ;
      RECT 0.0000 10.6780 59.8220 17.2100 ;
      RECT 0.0000 9.0780 58.9220 10.6780 ;
      RECT 0.0000 0.9000 59.8220 9.0780 ;
      RECT 0.0000 0.0000 22.8800 0.9000 ;
      RECT 35.4170 0.0000 59.8220 9.0780 ;
      RECT 35.4170 0.0000 59.8220 0.9000 ;
    LAYER M4 ;
      RECT 58.3210 225.3140 59.8220 226.8670 ;
      RECT 0.0000 200.8640 59.8220 206.5540 ;
      RECT 0.0000 192.0330 58.9250 206.5540 ;
      RECT 0.0000 181.6490 58.9230 206.5540 ;
      RECT 0.0000 199.2640 58.9250 200.8640 ;
      RECT 0.0000 197.7320 58.9380 199.2640 ;
      RECT 0.0000 192.0330 58.9380 199.2640 ;
      RECT 0.0000 192.0330 59.8220 197.7320 ;
      RECT 0.0000 190.4330 58.9230 192.0330 ;
      RECT 0.0000 188.8700 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 183.2150 59.8220 188.8700 ;
      RECT 0.0000 181.6490 58.9250 183.2150 ;
      RECT 0.0000 180.0490 58.9220 181.6490 ;
      RECT 0.0000 30.3170 59.8220 180.0490 ;
      RECT 0.0000 27.9920 58.9220 30.3170 ;
      RECT 0.0000 19.5650 59.8220 27.9920 ;
      RECT 0.0000 17.2100 58.9220 19.5650 ;
      RECT 0.0000 10.6780 59.8220 17.2100 ;
      RECT 0.0000 9.0780 58.9220 10.6780 ;
      RECT 0.0000 0.9000 59.8220 9.0780 ;
      RECT 0.0000 0.0000 22.8800 0.9000 ;
      RECT 35.4170 0.0000 59.8220 9.0780 ;
      RECT 35.4170 0.0000 59.8220 0.9000 ;
      RECT 0.0000 228.4670 59.8220 244.5640 ;
      RECT 0.0000 208.1540 58.9280 244.5640 ;
      RECT 0.0000 0.0000 22.8800 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 223.1530 58.9280 228.4670 ;
      RECT 0.0000 208.1540 59.8220 223.1530 ;
      RECT 0.0000 206.5540 58.9220 208.1540 ;
    LAYER M3 ;
      RECT 58.3210 225.3140 59.8220 226.8670 ;
      RECT 0.0000 200.8640 59.8220 206.5540 ;
      RECT 0.0000 192.0330 58.9250 206.5540 ;
      RECT 0.0000 181.6490 58.9230 206.5540 ;
      RECT 0.0000 199.2640 58.9250 200.8640 ;
      RECT 0.0000 197.7320 58.9380 199.2640 ;
      RECT 0.0000 192.0330 58.9380 199.2640 ;
      RECT 0.0000 192.0330 59.8220 197.7320 ;
      RECT 0.0000 190.4330 58.9230 192.0330 ;
      RECT 0.0000 188.8700 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 181.6490 58.9250 190.4330 ;
      RECT 0.0000 183.2150 59.8220 188.8700 ;
      RECT 0.0000 181.6490 58.9250 183.2150 ;
      RECT 0.0000 180.0490 58.9220 181.6490 ;
      RECT 0.0000 30.3170 59.8220 180.0490 ;
      RECT 0.0000 27.9920 58.9220 30.3170 ;
      RECT 0.0000 19.5650 59.8220 27.9920 ;
      RECT 0.0000 17.2100 58.9220 19.5650 ;
      RECT 0.0000 10.6780 59.8220 17.2100 ;
      RECT 0.0000 9.0780 58.9220 10.6780 ;
      RECT 0.0000 0.9000 59.8220 9.0780 ;
      RECT 0.0000 0.0000 22.8800 0.9000 ;
      RECT 35.4170 0.0000 59.8220 9.0780 ;
      RECT 35.4170 0.0000 59.8220 0.9000 ;
      RECT 0.0000 228.4670 59.8220 244.5640 ;
      RECT 0.0000 208.1540 58.9280 244.5640 ;
      RECT 0.0000 0.0000 22.8800 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 0.9000 58.9220 244.5640 ;
      RECT 0.0000 223.1530 58.9280 228.4670 ;
      RECT 0.0000 208.1540 59.8220 223.1530 ;
      RECT 0.0000 206.5540 58.9220 208.1540 ;
  END
END SRAMLP1RW512x8

MACRO SRAMLP1RW512x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 197.623 BY 258.787 ;
  SYMMETRY X Y R90 ;

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 175.3010 0.0000 175.5010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.3010 0.0000 175.5010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.3010 0.0000 175.5010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 175.3010 0.0000 175.5010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 175.3010 0.0000 175.5010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 41.0530 197.6230 41.2530 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 41.0530 197.6230 41.2530 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 41.0530 197.6230 41.2530 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 41.0530 197.6230 41.2530 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 41.0530 197.6230 41.2530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[8]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 16.9990 197.6230 17.1990 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 16.9990 197.6230 17.1990 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 16.9990 197.6230 17.1990 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 16.9990 197.6230 17.1990 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 16.9990 197.6230 17.1990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 16.4880 197.6230 16.6880 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 16.4880 197.6230 16.6880 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 16.4880 197.6230 16.6880 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 16.4880 197.6230 16.6880 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 16.4880 197.6230 16.6880 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 193.9170 258.4870 194.2160 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.4170 258.4870 0.7170 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3160 258.4870 1.6150 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.1170 258.4870 192.4160 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.0170 258.4870 193.3160 258.7870 ;
    END
  END VDD

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 133.5600 0.0000 133.7600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.5600 0.0000 133.7600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.5600 0.0000 133.7600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 133.5600 0.0000 133.7600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 133.5600 0.0000 133.7600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[0]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 134.2610 0.0000 134.4610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.2610 0.0000 134.4610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.2610 0.0000 134.4610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.2610 0.0000 134.4610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 134.2610 0.0000 134.4610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 134.9280 0.0000 135.1280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.9280 0.0000 135.1280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.9280 0.0000 135.1280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.9280 0.0000 135.1280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 134.9280 0.0000 135.1280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[1]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 135.6290 0.0000 135.8290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 135.6290 0.0000 135.8290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 135.6290 0.0000 135.8290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 135.6290 0.0000 135.8290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 135.6290 0.0000 135.8290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 136.2960 0.0000 136.4960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.2960 0.0000 136.4960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.2960 0.0000 136.4960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 136.2960 0.0000 136.4960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 136.2960 0.0000 136.4960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[2]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 136.9970 0.0000 137.1970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.9970 0.0000 137.1970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.9970 0.0000 137.1970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 136.9970 0.0000 137.1970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 136.9970 0.0000 137.1970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 137.6640 0.0000 137.8640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.6640 0.0000 137.8640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.6640 0.0000 137.8640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 137.6640 0.0000 137.8640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 137.6640 0.0000 137.8640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[3]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 138.3650 0.0000 138.5650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.3650 0.0000 138.5650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.3650 0.0000 138.5650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 138.3650 0.0000 138.5650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 138.3650 0.0000 138.5650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 139.0320 0.0000 139.2320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.0320 0.0000 139.2320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.0320 0.0000 139.2320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 139.0320 0.0000 139.2320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 139.0320 0.0000 139.2320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[4]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 139.7330 0.0000 139.9330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.7330 0.0000 139.9330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.7330 0.0000 139.9330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 139.7330 0.0000 139.9330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 139.7330 0.0000 139.9330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 140.4000 0.0000 140.6000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 140.4000 0.0000 140.6000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 140.4000 0.0000 140.6000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 140.4000 0.0000 140.6000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 140.4000 0.0000 140.6000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[5]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 141.1010 0.0000 141.3010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.1010 0.0000 141.3010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.1010 0.0000 141.3010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 141.1010 0.0000 141.3010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 141.1010 0.0000 141.3010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 141.7720 0.0000 141.9720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.7720 0.0000 141.9720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.7720 0.0000 141.9720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 141.7720 0.0000 141.9720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 141.7720 0.0000 141.9720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[6]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 142.4690 0.0000 142.6690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.4690 0.0000 142.6690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.4690 0.0000 142.6690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 142.4690 0.0000 142.6690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 142.4690 0.0000 142.6690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 172.5650 0.0000 172.7650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 172.5650 0.0000 172.7650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 172.5650 0.0000 172.7650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 172.5650 0.0000 172.7650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 172.5650 0.0000 172.7650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 9.7900 197.6230 9.9900 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 9.7930 197.6230 9.9930 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 9.7930 197.6230 9.9930 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 9.7930 197.6230 9.9930 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 9.7930 197.6230 9.9930 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 174.5980 0.0000 174.7980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 174.5980 0.0000 174.7980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 174.5980 0.0000 174.7980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 174.5980 0.0000 174.7980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 174.5980 0.0000 174.7980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[30]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 173.2340 0.0000 173.4340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.2340 0.0000 173.4340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.2350 0.0000 173.4350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 173.2350 0.0000 173.4350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 173.2350 0.0000 173.4350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[29]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 173.9330 0.0000 174.1330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.9330 0.0000 174.1330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.9330 0.0000 174.1330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 173.9330 0.0000 174.1330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 173.9330 0.0000 174.1330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 202.5220 197.6230 202.7220 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 202.5220 197.6230 202.7220 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 202.5220 197.6230 202.7220 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 202.5220 197.6230 202.7220 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 202.5220 197.6230 202.7220 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 204.1100 197.6230 204.3100 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 204.1100 197.6230 204.3100 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 204.1100 197.6230 204.3100 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 204.1100 197.6230 204.3100 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 204.1100 197.6230 204.3100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 211.3400 197.6230 211.5400 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 211.3400 197.6230 211.5400 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 211.3400 197.6230 211.5400 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 211.3400 197.6230 211.5400 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 211.3400 197.6230 211.5400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 212.9380 197.6230 213.1380 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 212.9380 197.6230 213.1380 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 212.9380 197.6230 213.1380 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 212.9380 197.6230 213.1380 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 212.9380 197.6230 213.1380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 220.1600 197.6230 220.3600 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 220.1600 197.6230 220.3600 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 220.1600 197.6230 220.3600 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 220.1600 197.6230 220.3600 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 220.1600 197.6230 220.3600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 176.6570 0.0000 176.8570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.6570 0.0000 176.8570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.6570 0.0000 176.8570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 176.6570 0.0000 176.8570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 176.6570 0.0000 176.8570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 195.2950 197.6230 195.4950 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 195.2950 197.6230 195.4950 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 195.2950 197.6230 195.4950 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 195.2950 197.6230 195.4950 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 195.2950 197.6230 195.4950 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2180 258.4870 2.5170 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.1170 258.4870 3.4180 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.3180 258.4870 190.6170 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.2180 258.4870 191.5180 258.7870 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 250.9220 197.6230 251.1220 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 250.9220 197.6230 251.1220 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 250.9220 197.6230 251.1220 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 250.9220 197.6230 251.1220 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 250.9220 197.6230 251.1220 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 247.7340 197.6230 247.9340 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 247.7340 197.6230 247.9340 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 247.7340 197.6230 247.9340 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 247.7340 197.6230 247.9340 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 247.7340 197.6230 247.9340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 247.2160 197.6230 247.4160 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 247.2160 197.6230 247.4160 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 247.2160 197.6230 247.4160 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 247.2160 197.6230 247.4160 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 247.2160 197.6230 247.4160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 193.7010 197.6230 193.9010 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 193.7010 197.6230 193.9010 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 193.7010 197.6230 193.9010 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 193.7010 197.6230 193.9010 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 193.7010 197.6230 193.9010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.4230 41.6140 197.6230 41.8140 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.4230 41.6140 197.6230 41.8140 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.4230 41.6140 197.6230 41.8140 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.4230 41.6140 197.6230 41.8140 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.4230 41.6140 197.6230 41.8140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.8930 0.0000 133.0930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.8930 0.0000 133.0930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.8930 0.0000 133.0930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.8930 0.0000 133.0930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.8930 0.0000 133.0930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 167.0930 0.0000 167.2930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.0930 0.0000 167.2930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.0930 0.0000 167.2930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 167.0930 0.0000 167.2930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 167.0930 0.0000 167.2930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 160.2530 0.0000 160.4530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.2530 0.0000 160.4530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.2530 0.0000 160.4530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 160.2530 0.0000 160.4530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 160.2530 0.0000 160.4530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 162.2870 0.0000 162.4870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 162.2870 0.0000 162.4870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 162.2870 0.0000 162.4870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 162.2870 0.0000 162.4870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 162.2870 0.0000 162.4870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[21]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 163.6580 0.0000 163.8580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 163.6580 0.0000 163.8580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 163.6600 0.0000 163.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 163.6600 0.0000 163.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 163.6600 0.0000 163.8600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[22]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 162.9890 0.0000 163.1890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 162.9890 0.0000 163.1890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 162.9890 0.0000 163.1890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 162.9890 0.0000 163.1890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 162.9890 0.0000 163.1890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 164.3570 0.0000 164.5570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.3570 0.0000 164.5570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.3570 0.0000 164.5570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 164.3570 0.0000 164.5570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 164.3570 0.0000 164.5570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 155.4470 0.0000 155.6470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 155.4470 0.0000 155.6470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 155.4470 0.0000 155.6470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 155.4470 0.0000 155.6470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 155.4470 0.0000 155.6470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[16]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 152.7120 0.0000 152.9120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.7120 0.0000 152.9120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.7120 0.0000 152.9120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 152.7120 0.0000 152.9120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 152.7120 0.0000 152.9120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[14]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 160.9190 0.0000 161.1190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.9190 0.0000 161.1190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.9190 0.0000 161.1190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 160.9190 0.0000 161.1190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 160.9190 0.0000 161.1190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[20]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 156.1490 0.0000 156.3490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.1490 0.0000 156.3490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.1490 0.0000 156.3490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 156.1490 0.0000 156.3490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 156.1490 0.0000 156.3490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 157.5170 0.0000 157.7170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 157.5170 0.0000 157.7170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 157.5170 0.0000 157.7170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 157.5170 0.0000 157.7170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 157.5170 0.0000 157.7170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 161.6210 0.0000 161.8210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.6210 0.0000 161.8210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.6210 0.0000 161.8210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 161.6210 0.0000 161.8210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 161.6210 0.0000 161.8210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.0780 0.0000 154.2780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.0780 0.0000 154.2780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.0780 0.0000 154.2780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.0780 0.0000 154.2780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.0780 0.0000 154.2780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[15]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 165.7250 0.0000 165.9250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.7250 0.0000 165.9250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.7250 0.0000 165.9250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 165.7250 0.0000 165.9250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 165.7250 0.0000 165.9250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 152.0450 0.0000 152.2450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.0450 0.0000 152.2450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.0450 0.0000 152.2450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 152.0450 0.0000 152.2450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 152.0450 0.0000 152.2450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 153.4130 0.0000 153.6130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.4130 0.0000 153.6130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.4130 0.0000 153.6130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 153.4130 0.0000 153.6130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 153.4130 0.0000 153.6130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.7810 0.0000 154.9810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.7810 0.0000 154.9810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.7810 0.0000 154.9810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.7810 0.0000 154.9810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.7810 0.0000 154.9810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 165.0260 0.0000 165.2260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.0260 0.0000 165.2260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.0260 0.0000 165.2260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 165.0260 0.0000 165.2260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 165.0260 0.0000 165.2260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[23]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 169.8290 0.0000 170.0290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.8290 0.0000 170.0290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.8290 0.0000 170.0290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 169.8290 0.0000 170.0290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 169.8290 0.0000 170.0290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 170.4950 0.0000 170.6950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 170.4950 0.0000 170.6950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 170.4950 0.0000 170.6950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 170.4950 0.0000 170.6950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 170.4950 0.0000 170.6950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[27]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 171.1970 0.0000 171.3970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.1970 0.0000 171.3970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.1970 0.0000 171.3970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 171.1970 0.0000 171.3970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 171.1970 0.0000 171.3970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 171.8640 0.0000 172.0640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.8640 0.0000 172.0640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.8640 0.0000 172.0640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 171.8640 0.0000 172.0640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 171.8640 0.0000 172.0640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[28]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 169.1270 0.0000 169.3270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.1270 0.0000 169.3270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.1270 0.0000 169.3270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 169.1270 0.0000 169.3270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 169.1270 0.0000 169.3270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[26]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 167.7590 0.0000 167.9590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.7590 0.0000 167.9590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.7590 0.0000 167.9590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 167.7590 0.0000 167.9590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 167.7590 0.0000 167.9590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[25]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.8850 0.0000 159.0850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.8850 0.0000 159.0850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.8850 0.0000 159.0850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 158.8850 0.0000 159.0850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 158.8850 0.0000 159.0850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 168.4610 0.0000 168.6610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.4610 0.0000 168.6610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.4610 0.0000 168.6610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 168.4610 0.0000 168.6610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 168.4610 0.0000 168.6610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 156.8160 0.0000 157.0160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.8160 0.0000 157.0160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.8160 0.0000 157.0160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 156.8160 0.0000 157.0160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 156.8160 0.0000 157.0160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[17]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 166.3920 0.0000 166.5920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 166.3920 0.0000 166.5920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 166.3920 0.0000 166.5920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 166.3920 0.0000 166.5920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 166.3920 0.0000 166.5920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[24]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 159.5550 0.0000 159.7550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 159.5550 0.0000 159.7550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 159.5550 0.0000 159.7550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 159.5550 0.0000 159.7550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 159.5550 0.0000 159.7550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[19]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.1840 0.0000 158.3840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.1840 0.0000 158.3840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.1840 0.0000 158.3840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 158.1840 0.0000 158.3840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 158.1840 0.0000 158.3840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[18]

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 1.7660 258.4870 2.0660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.8670 258.4870 1.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.5680 258.4870 3.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.6680 258.4870 2.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.4680 258.4870 4.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.3670 258.4870 5.6680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.0670 258.4870 8.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.1670 258.4870 7.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.2670 258.4870 6.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.9680 258.4870 9.2680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.7680 258.4870 11.0690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.6670 258.4870 11.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.8670 258.4870 10.1660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.5670 258.4870 12.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.2680 258.4870 15.5690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.9680 258.4870 18.2680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.4680 258.4870 13.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.3670 258.4870 14.6660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.1670 258.4870 16.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.0670 258.4870 17.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.5670 258.4870 21.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.4680 258.4870 22.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.6670 258.4870 20.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.7680 258.4870 20.0690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.8670 258.4870 19.1660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.8670 258.4870 28.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.9670 258.4870 27.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.1670 258.4870 25.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.2670 258.4870 24.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.3670 258.4870 23.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.0680 258.4870 26.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.3660 258.4870 32.6660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.4670 258.4870 31.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.5670 258.4870 30.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.7670 258.4870 29.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.6680 258.4870 29.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.1660 258.4870 34.4660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.2670 258.4870 33.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.8680 258.4870 37.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.9680 258.4870 36.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.0680 258.4870 35.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.7670 258.4870 38.0680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.3680 258.4870 41.6680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.4670 258.4870 40.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.5670 258.4870 39.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.2670 258.4870 42.5660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.6670 258.4870 38.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.8680 258.4870 46.1680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.7670 258.4870 47.0660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.1680 258.4870 43.4690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.0670 258.4870 44.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.9670 258.4870 45.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.2670 258.4870 51.5660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.6680 258.4870 47.9690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.3680 258.4870 50.6680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.5670 258.4870 48.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.4670 258.4870 49.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.6670 258.4870 56.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.7670 258.4870 56.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.9670 258.4870 54.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.8680 258.4870 55.1680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.0670 258.4870 53.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.1680 258.4870 52.4690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.1670 258.4870 61.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.2670 258.4870 60.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.3670 258.4870 59.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.5670 258.4870 57.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.4680 258.4870 58.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.7660 258.4870 65.0660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.8670 258.4870 64.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.9670 258.4870 63.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.6670 258.4870 65.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.0680 258.4870 62.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.5660 258.4870 66.8660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.2680 258.4870 69.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.1670 258.4870 70.4680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.3680 258.4870 68.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.4680 258.4870 67.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.0670 258.4870 71.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.7680 258.4870 74.0680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.5680 258.4870 75.8690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.8670 258.4870 73.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.9670 258.4870 72.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.6670 258.4870 74.9660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.0680 258.4870 80.3690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.2680 258.4870 78.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.1670 258.4870 79.4660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.4670 258.4870 76.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.3670 258.4870 77.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.4670 258.4870 85.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.5680 258.4870 84.8690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.6670 258.4870 83.9660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.7680 258.4870 83.0680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.9670 258.4870 81.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.8670 258.4870 82.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.1670 258.4870 88.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.3670 258.4870 86.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.2680 258.4870 87.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.9670 258.4870 90.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.0670 258.4870 89.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.4680 258.4870 94.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.8680 258.4870 91.1680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.5670 258.4870 93.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.6670 258.4870 92.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.7670 258.4870 92.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.0670 258.4870 98.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.9660 258.4870 99.2660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.1660 258.4870 97.4660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.2670 258.4870 96.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.3670 258.4870 95.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.8680 258.4870 100.1680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.6680 258.4870 101.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.5670 258.4870 102.8680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.3670 258.4870 104.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.7680 258.4870 101.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.4670 258.4870 103.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.1680 258.4870 106.4680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.9680 258.4870 108.2690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.8670 258.4870 109.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.2670 258.4870 105.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.0670 258.4870 107.3660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.7670 258.4870 110.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.4680 258.4870 112.7690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.5670 258.4870 111.8660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.3670 258.4870 113.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.2670 258.4870 114.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.6680 258.4870 110.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.8670 258.4870 118.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.9680 258.4870 117.2690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.0670 258.4870 116.3660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.1680 258.4870 115.4680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.7670 258.4870 119.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.2680 258.4870 123.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.6680 258.4870 119.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.1670 258.4870 124.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.3670 258.4870 122.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.4670 258.4870 121.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.5670 258.4870 120.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.8680 258.4870 127.1680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.6670 258.4870 128.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.7670 258.4870 128.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.9670 258.4870 126.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.0670 258.4870 125.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.4670 258.4870 130.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.3660 258.4870 131.6660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.5660 258.4870 129.8660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.1680 258.4870 133.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.2680 258.4870 132.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.0680 258.4870 134.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.9670 258.4870 135.2680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.5680 258.4870 138.8680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.6670 258.4870 137.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.7670 258.4870 137.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.8670 258.4870 136.1680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.3680 258.4870 140.6690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.2670 258.4870 141.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.4670 258.4870 139.7660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.1670 258.4870 142.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.0680 258.4870 143.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.8680 258.4870 145.1690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.5680 258.4870 147.8680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.9670 258.4870 144.2660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.7670 258.4870 146.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.6670 258.4870 146.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.0680 258.4870 152.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.2670 258.4870 150.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.3680 258.4870 149.6690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.4670 258.4870 148.7660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.9670 258.4870 153.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.1670 258.4870 151.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.6680 258.4870 155.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.4670 258.4870 157.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.5670 258.4870 156.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.7670 258.4870 155.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.8670 258.4870 154.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.2680 258.4870 159.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.9660 258.4870 162.2660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.0670 258.4870 161.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.1670 258.4870 160.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.3670 258.4870 158.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.8670 258.4870 163.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.4680 258.4870 166.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.3670 258.4870 167.6680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 163.7660 258.4870 164.0660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.5680 258.4870 165.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.6680 258.4870 164.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.9680 258.4870 171.2680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.0670 258.4870 170.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.1670 258.4870 169.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.8670 258.4870 172.1660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.2670 258.4870 168.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.3670 258.4870 176.6660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.7680 258.4870 173.0690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.6670 258.4870 173.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 174.5670 258.4870 174.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.4680 258.4870 175.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.7680 258.4870 182.0690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.8670 258.4870 181.1660 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.2680 258.4870 177.5690 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.9680 258.4870 180.2680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.1670 258.4870 178.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.0670 258.4870 179.3670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.4680 258.4870 184.7680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.6670 258.4870 182.9670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.2670 258.4870 186.5670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 185.3670 258.4870 185.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.5670 258.4870 183.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.0680 258.4870 188.3680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.7670 258.4870 191.0670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.8670 258.4870 190.1670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.9670 258.4870 189.2670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.5670 258.4870 192.8670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.4670 258.4870 193.7670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.3670 258.4870 194.6670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.1670 258.4870 196.4670 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.6680 258.4870 191.9680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 195.2680 258.4870 195.5680 258.7870 ;
    END
    PORT
      LAYER M5 ;
        RECT 187.1670 258.4870 187.4670 258.7870 ;
    END
  END VSS

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 143.1370 0.0000 143.3370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.1370 0.0000 143.3370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.1370 0.0000 143.3370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 143.1370 0.0000 143.3370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 143.1370 0.0000 143.3370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[7]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 143.8370 0.0000 144.0370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.8370 0.0000 144.0370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.8370 0.0000 144.0370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 143.8370 0.0000 144.0370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 143.8370 0.0000 144.0370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 144.5110 0.0000 144.7110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.5110 0.0000 144.7110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.5110 0.0000 144.7110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 144.5110 0.0000 144.7110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 144.5110 0.0000 144.7110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[8]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 145.2050 0.0000 145.4050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.2050 0.0000 145.4050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.2050 0.0000 145.4050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 145.2050 0.0000 145.4050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 145.2050 0.0000 145.4050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 145.8790 0.0000 146.0790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.8790 0.0000 146.0790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.8790 0.0000 146.0790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 145.8790 0.0000 146.0790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 145.8790 0.0000 146.0790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[9]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 146.5730 0.0000 146.7730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.5730 0.0000 146.7730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.5730 0.0000 146.7730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 146.5730 0.0000 146.7730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 146.5730 0.0000 146.7730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 147.2400 0.0000 147.4400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.2400 0.0000 147.4400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.2400 0.0000 147.4400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 147.2400 0.0000 147.4400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 147.2400 0.0000 147.4400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[10]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 147.9410 0.0000 148.1410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.9410 0.0000 148.1410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.9410 0.0000 148.1410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 147.9410 0.0000 148.1410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 147.9410 0.0000 148.1410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.6080 0.0000 148.8080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.6080 0.0000 148.8080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.6080 0.0000 148.8080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.6080 0.0000 148.8080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.6080 0.0000 148.8080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[11]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 149.3090 0.0000 149.5090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.3090 0.0000 149.5090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.3090 0.0000 149.5090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 149.3090 0.0000 149.5090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 149.9760 0.0000 150.1760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.9760 0.0000 150.1760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.9760 0.0000 150.1760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 149.9760 0.0000 150.1760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 149.9760 0.0000 150.1760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[12]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.6770 0.0000 150.8770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.6770 0.0000 150.8770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.6770 0.0000 150.8770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.6770 0.0000 150.8770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.6770 0.0000 150.8770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 151.3420 0.0000 151.5420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 151.3420 0.0000 151.5420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 151.3420 0.0000 151.5420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 151.3420 0.0000 151.5420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 151.3420 0.0000 151.5420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[13]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 175.9720 0.0000 176.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.9720 0.0000 176.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.9720 0.0000 176.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 175.9720 0.0000 176.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 175.9720 0.0000 176.1720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[31]
  OBS
    LAYER M1 ;
      RECT 196.8230 203.3220 197.6230 203.5100 ;
      RECT 196.8230 212.1400 197.6230 212.3380 ;
      RECT 196.1220 248.5340 197.6230 250.3220 ;
      RECT 0.0000 251.7220 197.6230 258.7870 ;
      RECT 0.0000 0.0000 132.2930 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 0.8000 196.8230 258.7870 ;
      RECT 0.0000 246.6160 196.8230 251.7220 ;
      RECT 0.0000 220.9600 197.6230 246.6160 ;
      RECT 0.0000 219.5600 196.8230 220.9600 ;
      RECT 0.0000 213.7380 197.6230 219.5600 ;
      RECT 0.0000 210.7400 196.8230 213.7380 ;
      RECT 0.0000 204.9100 197.6230 210.7400 ;
      RECT 0.0000 201.9220 196.8230 204.9100 ;
      RECT 0.0000 196.0950 197.6230 201.9220 ;
      RECT 0.0000 193.1010 196.8230 196.0950 ;
      RECT 0.0000 42.4140 197.6230 193.1010 ;
      RECT 0.0000 40.4530 196.8230 42.4140 ;
      RECT 0.0000 17.7990 197.6230 40.4530 ;
      RECT 0.0000 15.8880 196.8230 17.7990 ;
      RECT 0.0000 10.5930 197.6230 15.8880 ;
      RECT 0.0000 9.1930 196.8230 10.5930 ;
      RECT 0.0000 0.8000 197.6230 9.1930 ;
      RECT 0.0000 0.0000 132.2930 0.8000 ;
      RECT 177.4570 0.0000 197.6230 9.1930 ;
      RECT 177.4570 0.0000 197.6230 0.8000 ;
      RECT 196.8230 194.5010 197.6230 194.6950 ;
    LAYER PO ;
      RECT 0.0000 0.0000 197.6230 258.7870 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 197.6230 258.7870 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 197.6230 258.7870 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 197.6230 258.7870 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 197.6230 258.7870 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 197.6230 258.7870 ;
    LAYER M5 ;
      RECT 197.1670 257.7870 197.6230 258.7870 ;
      RECT 196.1220 248.6340 197.6230 250.2220 ;
      RECT 0.0000 251.8220 197.6230 257.7870 ;
      RECT 0.0000 0.0000 132.1930 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 0.9000 196.7230 257.7870 ;
      RECT 0.0000 246.5160 196.7230 251.8220 ;
      RECT 0.0000 221.0600 197.6230 246.5160 ;
      RECT 0.0000 219.4600 196.7230 221.0600 ;
      RECT 0.0000 213.8380 197.6230 219.4600 ;
      RECT 0.0000 210.6400 196.7230 213.8380 ;
      RECT 0.0000 205.0100 197.6230 210.6400 ;
      RECT 0.0000 201.8220 196.7230 205.0100 ;
      RECT 0.0000 196.1950 197.6230 201.8220 ;
      RECT 0.0000 193.0010 196.7230 196.1950 ;
      RECT 0.0000 42.5140 197.6230 193.0010 ;
      RECT 0.0000 40.3530 196.7230 42.5140 ;
      RECT 0.0000 17.8990 197.6230 40.3530 ;
      RECT 0.0000 15.7880 196.7230 17.8990 ;
      RECT 0.0000 10.6900 197.6230 15.7880 ;
      RECT 0.0000 9.0900 196.7230 10.6900 ;
      RECT 0.0000 0.9000 197.6230 9.0900 ;
      RECT 0.0000 0.0000 132.1930 0.9000 ;
      RECT 177.5570 0.0000 197.6230 9.0900 ;
      RECT 177.5570 0.0000 197.6230 0.9000 ;
    LAYER M4 ;
      RECT 196.1220 248.6340 197.6230 250.2220 ;
      RECT 0.0000 251.8220 197.6230 258.7870 ;
      RECT 0.0000 0.0000 132.1930 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 246.5160 196.7230 251.8220 ;
      RECT 0.0000 221.0600 197.6230 246.5160 ;
      RECT 0.0000 219.4600 196.7230 221.0600 ;
      RECT 0.0000 213.8380 197.6230 219.4600 ;
      RECT 0.0000 210.6400 196.7230 213.8380 ;
      RECT 0.0000 205.0100 197.6230 210.6400 ;
      RECT 0.0000 201.8220 196.7230 205.0100 ;
      RECT 0.0000 196.1950 197.6230 201.8220 ;
      RECT 0.0000 193.0010 196.7230 196.1950 ;
      RECT 0.0000 42.5140 197.6230 193.0010 ;
      RECT 0.0000 40.3530 196.7230 42.5140 ;
      RECT 0.0000 17.8990 197.6230 40.3530 ;
      RECT 0.0000 15.7880 196.7230 17.8990 ;
      RECT 0.0000 10.6930 197.6230 15.7880 ;
      RECT 0.0000 9.0930 196.7230 10.6930 ;
      RECT 0.0000 0.9000 197.6230 9.0930 ;
      RECT 0.0000 0.0000 132.1930 0.9000 ;
      RECT 177.5570 0.0000 197.6230 9.0930 ;
      RECT 177.5570 0.0000 197.6230 0.9000 ;
    LAYER M3 ;
      RECT 196.1220 248.6340 197.6230 250.2220 ;
      RECT 0.0000 251.8220 197.6230 258.7870 ;
      RECT 0.0000 0.0000 132.1930 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 246.5160 196.7230 251.8220 ;
      RECT 0.0000 221.0600 197.6230 246.5160 ;
      RECT 0.0000 219.4600 196.7230 221.0600 ;
      RECT 0.0000 213.8380 197.6230 219.4600 ;
      RECT 0.0000 210.6400 196.7230 213.8380 ;
      RECT 0.0000 205.0100 197.6230 210.6400 ;
      RECT 0.0000 201.8220 196.7230 205.0100 ;
      RECT 0.0000 196.1950 197.6230 201.8220 ;
      RECT 0.0000 193.0010 196.7230 196.1950 ;
      RECT 0.0000 42.5140 197.6230 193.0010 ;
      RECT 0.0000 40.3530 196.7230 42.5140 ;
      RECT 0.0000 17.8990 197.6230 40.3530 ;
      RECT 0.0000 15.7880 196.7230 17.8990 ;
      RECT 0.0000 10.6930 197.6230 15.7880 ;
      RECT 0.0000 9.0930 196.7230 10.6930 ;
      RECT 0.0000 0.9000 197.6230 9.0930 ;
      RECT 0.0000 0.0000 132.1930 0.9000 ;
      RECT 177.5570 0.0000 197.6230 9.0930 ;
      RECT 177.5570 0.0000 197.6230 0.9000 ;
    LAYER M2 ;
      RECT 196.1220 248.6340 197.6230 250.2220 ;
      RECT 0.0000 251.8220 197.6230 258.7870 ;
      RECT 0.0000 0.0000 132.1930 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 0.9000 196.7230 258.7870 ;
      RECT 0.0000 246.5160 196.7230 251.8220 ;
      RECT 0.0000 221.0600 197.6230 246.5160 ;
      RECT 0.0000 219.4600 196.7230 221.0600 ;
      RECT 0.0000 213.8380 197.6230 219.4600 ;
      RECT 0.0000 210.6400 196.7230 213.8380 ;
      RECT 0.0000 205.0100 197.6230 210.6400 ;
      RECT 0.0000 201.8220 196.7230 205.0100 ;
      RECT 0.0000 196.1950 197.6230 201.8220 ;
      RECT 0.0000 193.0010 196.7230 196.1950 ;
      RECT 0.0000 42.5140 197.6230 193.0010 ;
      RECT 0.0000 40.3530 196.7230 42.5140 ;
      RECT 0.0000 17.8990 197.6230 40.3530 ;
      RECT 0.0000 15.7880 196.7230 17.8990 ;
      RECT 0.0000 10.6930 197.6230 15.7880 ;
      RECT 0.0000 9.0930 196.7230 10.6930 ;
      RECT 0.0000 0.9000 197.6230 9.0930 ;
      RECT 0.0000 0.0000 132.1930 0.9000 ;
      RECT 177.5570 0.0000 197.6230 9.0930 ;
      RECT 177.5570 0.0000 197.6230 0.9000 ;
  END
END SRAMLP1RW512x32

MACRO SRAMLP1RW512x128
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 723.182 BY 309.594 ;
  SYMMETRY X Y R90 ;

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 539.1290 0.0000 539.3290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 539.1290 0.0000 539.3290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 539.1290 0.0000 539.3290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 539.1290 0.0000 539.3290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 539.1290 0.0000 539.3290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 539.8140 0.0000 540.0140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 539.8140 0.0000 540.0140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 539.8140 0.0000 540.0140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 539.8140 0.0000 540.0140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 539.8140 0.0000 540.0140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[9]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 537.7610 0.0000 537.9610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 537.7610 0.0000 537.9610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 537.7610 0.0000 537.9610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 537.7610 0.0000 537.9610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 537.7610 0.0000 537.9610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 538.4460 0.0000 538.6460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 538.4460 0.0000 538.6460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 538.4460 0.0000 538.6460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 538.4460 0.0000 538.6460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 538.4460 0.0000 538.6460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[8]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 537.0780 0.0000 537.2780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 537.0780 0.0000 537.2780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 537.0780 0.0000 537.2780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 537.0780 0.0000 537.2780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 537.0780 0.0000 537.2780 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[7]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 542.5500 0.0000 542.7500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 542.5500 0.0000 542.7500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 542.5500 0.0000 542.7500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 542.5500 0.0000 542.7500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 542.5500 0.0000 542.7500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[11]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 547.3370 0.0000 547.5370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 547.3370 0.0000 547.5370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 547.3370 0.0000 547.5370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 547.3370 0.0000 547.5370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 547.3370 0.0000 547.5370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 548.0220 0.0000 548.2220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 548.0220 0.0000 548.2220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 548.0220 0.0000 548.2220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 548.0220 0.0000 548.2220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 548.0220 0.0000 548.2220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[15]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 545.9690 0.0000 546.1690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 545.9690 0.0000 546.1690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 545.9690 0.0000 546.1690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 545.9690 0.0000 546.1690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 545.9690 0.0000 546.1690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 546.6540 0.0000 546.8540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 546.6540 0.0000 546.8540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 546.6540 0.0000 546.8540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 546.6540 0.0000 546.8540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 546.6540 0.0000 546.8540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[14]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 545.2860 0.0000 545.4860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 545.2860 0.0000 545.4860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 545.2860 0.0000 545.4860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 545.2860 0.0000 545.4860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 545.2860 0.0000 545.4860 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[13]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 543.9180 0.0000 544.1180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 543.9180 0.0000 544.1180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 543.9180 0.0000 544.1180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 543.9180 0.0000 544.1180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 543.9180 0.0000 544.1180 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[12]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 544.6010 0.0000 544.8010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 544.6010 0.0000 544.8010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 544.6010 0.0000 544.8010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 544.6010 0.0000 544.8010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 544.6010 0.0000 544.8010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 543.2330 0.0000 543.4330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 543.2330 0.0000 543.4330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 543.2330 0.0000 543.4330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 543.2330 0.0000 543.4330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 543.2330 0.0000 543.4330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 550.7580 0.0000 550.9580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 550.7580 0.0000 550.9580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 550.7580 0.0000 550.9580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 550.7580 0.0000 550.9580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 550.7580 0.0000 550.9580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[17]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9880 288.3990 723.1820 288.5990 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9880 288.3990 723.1820 288.5990 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9880 288.3990 723.1820 288.5990 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9880 288.3990 723.1820 288.5990 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9880 288.3990 723.1820 288.5990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9880 291.6510 723.1820 291.8510 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9880 291.6510 723.1820 291.8510 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9880 291.6510 723.1820 291.8510 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9880 291.6510 723.1820 291.8510 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9880 291.6510 723.1820 291.8510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 17.2900 723.1820 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 17.2900 723.1820 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 17.2900 723.1820 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 17.2900 723.1820 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 17.2900 723.1820 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 708.2990 309.2940 708.5990 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 709.1990 309.2940 709.4990 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 710.1000 309.2940 710.4000 309.5940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 529.5530 0.0000 529.7530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 529.5530 0.0000 529.7530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 529.5530 0.0000 529.7530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 529.5530 0.0000 529.7530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 529.5530 0.0000 529.7530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 530.2380 0.0000 530.4380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 530.2380 0.0000 530.4380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 530.2380 0.0000 530.4380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 530.2380 0.0000 530.4380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 530.2380 0.0000 530.4380 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[2]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 527.5020 0.0000 527.7020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 527.5020 0.0000 527.7020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 527.5020 0.0000 527.7020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 527.5020 0.0000 527.7020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 527.5020 0.0000 527.7020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[0]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 528.8700 0.0000 529.0700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 528.8700 0.0000 529.0700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 528.8700 0.0000 529.0700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 528.8700 0.0000 529.0700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 528.8700 0.0000 529.0700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[1]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 528.1850 0.0010 528.3850 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 528.1850 0.0010 528.3850 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 528.1850 0.0000 528.3850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 528.1850 0.0000 528.3850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 528.1850 0.0000 528.3850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 526.8170 0.0000 527.0170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 526.8170 0.0000 527.0170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 526.8170 0.0000 527.0170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 526.8170 0.0000 527.0170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 526.8170 0.0000 527.0170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 532.9740 0.0000 533.1740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 532.9740 0.0000 533.1740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 532.9740 0.0000 533.1740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 532.9740 0.0000 533.1740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 532.9740 0.0000 533.1740 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[4]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 532.2890 0.0000 532.4890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 532.2890 0.0000 532.4890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 532.2890 0.0000 532.4890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 532.2890 0.0000 532.4890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 532.2890 0.0000 532.4890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 531.6060 0.0000 531.8060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 531.6060 0.0000 531.8060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 531.6060 0.0000 531.8060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 531.6060 0.0000 531.8060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 531.6060 0.0000 531.8060 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[3]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 530.9210 0.0000 531.1210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 530.9210 0.0000 531.1210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 530.9210 0.0000 531.1210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 530.9210 0.0000 531.1210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 530.9210 0.0000 531.1210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 535.7100 0.0000 535.9100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 535.7100 0.0000 535.9100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 535.7100 0.0000 535.9100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 535.7100 0.0000 535.9100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 535.7100 0.0000 535.9100 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[6]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 535.0250 0.0000 535.2250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 535.0250 0.0000 535.2250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 535.0250 0.0000 535.2250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 535.0250 0.0000 535.2250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 535.0250 0.0000 535.2250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 534.3420 0.0000 534.5420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 534.3420 0.0000 534.5420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 534.3420 0.0000 534.5420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 534.3420 0.0000 534.5420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 534.3420 0.0000 534.5420 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[5]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 533.6570 0.0000 533.8570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 533.6570 0.0000 533.8570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 533.6570 0.0000 533.8570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 533.6570 0.0000 533.8570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 533.6570 0.0000 533.8570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 245.5700 723.1820 245.7700 ;
    END
    PORT
      LAYER M5 ;
        RECT 722.9820 247.1600 723.1820 247.3600 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 247.1600 723.1820 247.3600 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 247.1600 723.1820 247.3600 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 247.1600 723.1820 247.3600 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 247.1600 723.1820 247.3600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 263.2060 723.1820 263.4060 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 263.2060 723.1820 263.4060 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 263.2060 723.1820 263.4060 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 263.2060 723.1820 263.4060 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 263.2060 723.1820 263.4060 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 255.9760 723.1820 256.1760 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 255.9760 723.1820 256.1760 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 255.9760 723.1820 256.1760 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 255.9760 723.1820 256.1760 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 255.9760 723.1820 256.1760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 264.7960 723.1820 264.9960 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 264.7960 723.1820 264.9960 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 264.7960 723.1820 264.9960 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 264.7960 723.1820 264.9960 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 264.7960 723.1820 264.9960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 254.3860 723.1820 254.5860 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 254.3860 723.1820 254.5860 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 254.3860 723.1820 254.5860 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 254.3860 723.1820 254.5860 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 254.3860 723.1820 254.5860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 272.0260 723.1820 272.2260 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 272.0260 723.1820 272.2260 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 272.0260 723.1820 272.2260 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 272.0260 723.1820 272.2260 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 272.0260 723.1820 272.2260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 719.1000 309.2940 719.4010 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 718.2000 309.2940 718.4990 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 717.2990 309.2940 717.5990 309.5940 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 3.1490 309.2940 3.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3500 309.2940 1.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.4500 309.2940 0.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2500 309.2940 2.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.0490 309.2940 4.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9490 309.2940 5.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.5500 309.2940 8.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.6490 309.2940 7.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.7500 309.2940 7.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8490 309.2940 6.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.4490 309.2940 9.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1490 309.2940 12.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.2500 309.2940 11.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.0500 309.2940 13.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.3490 309.2940 10.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.5500 309.2940 17.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.6500 309.2940 16.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.9490 309.2940 14.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4500 309.2940 18.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.8490 309.2940 15.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.7500 309.2940 16.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.1490 309.2940 21.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.3490 309.2940 19.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.9500 309.2940 23.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.0490 309.2940 22.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.2490 309.2940 20.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.6490 309.2940 25.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.7500 309.2940 25.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.8490 309.2940 24.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.4500 309.2940 27.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.5490 309.2940 26.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.8500 309.2940 33.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.3490 309.2940 28.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.2500 309.2940 29.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.1490 309.2940 30.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.0490 309.2940 31.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.9500 309.2940 32.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.3490 309.2940 37.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.5490 309.2940 35.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.7500 309.2940 34.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.6500 309.2940 34.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.4490 309.2940 36.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.8490 309.2940 42.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.9500 309.2940 41.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.0490 309.2940 40.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.1500 309.2940 39.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.2490 309.2940 38.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.5490 309.2940 44.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.6500 309.2940 43.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.4500 309.2940 45.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.3490 309.2940 46.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.7490 309.2940 43.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.2490 309.2940 47.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.7490 309.2940 52.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.9500 309.2940 50.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.0500 309.2940 49.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.8500 309.2940 51.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.1500 309.2940 48.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.5490 309.2940 53.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.2490 309.2940 56.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.3500 309.2940 55.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.4490 309.2940 54.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.6490 309.2940 52.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.0490 309.2940 58.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.1500 309.2940 57.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.7490 309.2940 61.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.8500 309.2940 60.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.6500 309.2940 61.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.9490 309.2940 59.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.1500 309.2940 66.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.2500 309.2940 65.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.5490 309.2940 62.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.4490 309.2940 63.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.3500 309.2940 64.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.7490 309.2940 70.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.9490 309.2940 68.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.0500 309.2940 67.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.8490 309.2940 69.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.6490 309.2940 70.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.2490 309.2940 74.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.3500 309.2940 73.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.4490 309.2940 72.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.0500 309.2940 76.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.5500 309.2940 71.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.1490 309.2940 75.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.9490 309.2940 77.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.8500 309.2940 78.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.7490 309.2940 79.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.6490 309.2940 79.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.5500 309.2940 80.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.1490 309.2940 84.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.3500 309.2940 82.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.4500 309.2940 81.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.2500 309.2940 83.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.0490 309.2940 85.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.9490 309.2940 86.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.4490 309.2940 90.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.5500 309.2940 89.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.6490 309.2940 88.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.7500 309.2940 88.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.8490 309.2940 87.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.1490 309.2940 93.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.2500 309.2940 92.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.0500 309.2940 94.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.9490 309.2940 95.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.3490 309.2940 91.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.3490 309.2940 100.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.5500 309.2940 98.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.6500 309.2940 97.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.4500 309.2940 99.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.8490 309.2940 96.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.7500 309.2940 97.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.1490 309.2940 102.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.8490 309.2940 105.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.9500 309.2940 104.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.2490 309.2940 101.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.0490 309.2940 103.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.6490 309.2940 106.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.7500 309.2940 106.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.3490 309.2940 109.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.4500 309.2940 108.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.5490 309.2940 107.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.7500 309.2940 115.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.8500 309.2940 114.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.2500 309.2940 110.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.1490 309.2940 111.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.0490 309.2940 112.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.9500 309.2940 113.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.3490 309.2940 118.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.5490 309.2940 116.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.6500 309.2940 115.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.4490 309.2940 117.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.2490 309.2940 119.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.8490 309.2940 123.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.9500 309.2940 122.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.0490 309.2940 121.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.1500 309.2940 120.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.7490 309.2940 124.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.5490 309.2940 125.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.6500 309.2940 124.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.4500 309.2940 126.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.3490 309.2940 127.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.2490 309.2940 128.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.1500 309.2940 129.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.7490 309.2940 133.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.9500 309.2940 131.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.0500 309.2940 130.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.8500 309.2940 132.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.6490 309.2940 133.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.5490 309.2940 134.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.1500 309.2940 138.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.2490 309.2940 137.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.3500 309.2940 136.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.4490 309.2940 135.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.0490 309.2940 139.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.7490 309.2940 142.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.8500 309.2940 141.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.6500 309.2940 142.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.5490 309.2940 143.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.9490 309.2940 140.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.1500 309.2940 147.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.2500 309.2940 146.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.0500 309.2940 148.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.4490 309.2940 144.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.3500 309.2940 145.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.7490 309.2940 151.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.9490 309.2940 149.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.5500 309.2940 152.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.8490 309.2940 150.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.6490 309.2940 151.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.2490 309.2940 155.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.3500 309.2940 154.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.9490 309.2940 158.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.4490 309.2940 153.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.0500 309.2940 157.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.1490 309.2940 156.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.4500 309.2940 162.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.8500 309.2940 159.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.7490 309.2940 160.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.6490 309.2940 160.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.5500 309.2940 161.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.9490 309.2940 167.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.1490 309.2940 165.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 163.3500 309.2940 163.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.2500 309.2940 164.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.0490 309.2940 166.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.4490 309.2940 171.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.5500 309.2940 170.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.6490 309.2940 169.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.7500 309.2940 169.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.3490 309.2940 172.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.8490 309.2940 168.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 174.1490 309.2940 174.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.2500 309.2940 173.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.0500 309.2940 175.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.9490 309.2940 176.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.8490 309.2940 177.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.3490 309.2940 181.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.5500 309.2940 179.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.6500 309.2940 178.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.4500 309.2940 180.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.7500 309.2940 178.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.2490 309.2940 182.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.1490 309.2940 183.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.7500 309.2940 187.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 185.8490 309.2940 186.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.9500 309.2940 185.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.0490 309.2940 184.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 187.6490 309.2940 187.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.3490 309.2940 190.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.4500 309.2940 189.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.2500 309.2940 191.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.5490 309.2940 188.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 195.7500 309.2940 196.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.8500 309.2940 195.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.1490 309.2940 192.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.6500 309.2940 196.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.0490 309.2940 193.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.9500 309.2940 194.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 199.3490 309.2940 199.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.5490 309.2940 197.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 201.1500 309.2940 201.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 198.4490 309.2940 198.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 200.2490 309.2940 200.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.8490 309.2940 204.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 202.9500 309.2940 203.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 202.0490 309.2940 202.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.6500 309.2940 205.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.7490 309.2940 205.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.0500 309.2940 211.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 206.5490 309.2940 206.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.4500 309.2940 207.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 208.3490 309.2940 208.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 209.2490 309.2940 209.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 210.1500 309.2940 210.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.5490 309.2940 215.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 213.7490 309.2940 214.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.9500 309.2940 212.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.8500 309.2940 213.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 214.6490 309.2940 214.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.0490 309.2940 220.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.1500 309.2940 219.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 218.2490 309.2940 218.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 217.3500 309.2940 217.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.4490 309.2940 216.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.7490 309.2940 223.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 221.8500 309.2940 222.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 223.6500 309.2940 223.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 224.5490 309.2940 224.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.9490 309.2940 221.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 225.4490 309.2940 225.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 229.9490 309.2940 230.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.1500 309.2940 228.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 227.2500 309.2940 227.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 229.0500 309.2940 229.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.3500 309.2940 226.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 231.7490 309.2940 232.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.4490 309.2940 234.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.5500 309.2940 233.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.8490 309.2940 231.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 232.6490 309.2940 232.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 236.2490 309.2940 236.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 235.3500 309.2940 235.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 238.9490 309.2940 239.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 238.0500 309.2940 238.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 239.8500 309.2940 240.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 237.1490 309.2940 237.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 244.3500 309.2940 244.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 243.4500 309.2940 243.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 240.7490 309.2940 241.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.6490 309.2940 241.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 242.5500 309.2940 242.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 247.9490 309.2940 248.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 246.1490 309.2940 246.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 245.2500 309.2940 245.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 247.0490 309.2940 247.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.8490 309.2940 249.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 252.4490 309.2940 252.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 251.5500 309.2940 251.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 250.6490 309.2940 250.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 254.2500 309.2940 254.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 249.7500 309.2940 250.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 253.3490 309.2940 253.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.1490 309.2940 255.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 256.0500 309.2940 256.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 256.9490 309.2940 257.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 257.8490 309.2940 258.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 258.7500 309.2940 259.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 262.3490 309.2940 262.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.5500 309.2940 260.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 259.6500 309.2940 259.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 261.4500 309.2940 261.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 263.2490 309.2940 263.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 264.1490 309.2940 264.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 268.6490 309.2940 268.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 267.7500 309.2940 268.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 266.8490 309.2940 267.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 265.9500 309.2940 266.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 265.0490 309.2940 265.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 271.3490 309.2940 271.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 270.4500 309.2940 270.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 272.2500 309.2940 272.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 273.1490 309.2940 273.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 269.5490 309.2940 269.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.5490 309.2940 278.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 276.7500 309.2940 277.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 275.8500 309.2940 276.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 277.6500 309.2940 277.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 274.0490 309.2940 274.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 274.9500 309.2940 275.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 280.3490 309.2940 280.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 283.0490 309.2940 283.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 282.1500 309.2940 282.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 279.4490 309.2940 279.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 281.2490 309.2940 281.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 284.8490 309.2940 285.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 283.9500 309.2940 284.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 287.5490 309.2940 287.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 286.6500 309.2940 286.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 285.7490 309.2940 286.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 292.9500 309.2940 293.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 292.0500 309.2940 292.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 288.4500 309.2940 288.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 289.3490 309.2940 289.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 290.2490 309.2940 290.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 291.1500 309.2940 291.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 296.5490 309.2940 296.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 294.7490 309.2940 295.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 293.8500 309.2940 294.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 295.6490 309.2940 295.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 297.4490 309.2940 297.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 301.0490 309.2940 301.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 300.1500 309.2940 300.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 299.2490 309.2940 299.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 298.3500 309.2940 298.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 301.9490 309.2940 302.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 303.7490 309.2940 304.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 302.8500 309.2940 303.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 304.6500 309.2940 304.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 305.5490 309.2940 305.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 306.4490 309.2940 306.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 307.3500 309.2940 307.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.9490 309.2940 311.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 309.1500 309.2940 309.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 308.2500 309.2940 308.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 310.0500 309.2940 310.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 311.8490 309.2940 312.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 312.7490 309.2940 313.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 316.3500 309.2940 316.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 315.4490 309.2940 315.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 314.5500 309.2940 314.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 313.6490 309.2940 313.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 317.2490 309.2940 317.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 319.9490 309.2940 320.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 319.0500 309.2940 319.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 320.8500 309.2940 321.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 321.7490 309.2940 322.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 318.1490 309.2940 318.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 325.3500 309.2940 325.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 324.4500 309.2940 324.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 326.2500 309.2940 326.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 322.6490 309.2940 322.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 323.5500 309.2940 323.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 327.1490 309.2940 327.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 328.9490 309.2940 329.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 330.7500 309.2940 331.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 328.0490 309.2940 328.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 329.8490 309.2940 330.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 333.4490 309.2940 333.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 332.5500 309.2940 332.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 336.1490 309.2940 336.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 331.6490 309.2940 331.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 335.2500 309.2940 335.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 334.3490 309.2940 334.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 340.6500 309.2940 340.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 337.0500 309.2940 337.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 337.9490 309.2940 338.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 338.8490 309.2940 339.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 339.7500 309.2940 340.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 343.3490 309.2940 343.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 341.5500 309.2940 341.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 345.1490 309.2940 345.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 342.4500 309.2940 342.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 344.2490 309.2940 344.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 349.6490 309.2940 349.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 348.7500 309.2940 349.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 347.8490 309.2940 348.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 346.9500 309.2940 347.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 350.5490 309.2940 350.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 346.0490 309.2940 346.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 352.3490 309.2940 352.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 351.4500 309.2940 351.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 353.2500 309.2940 353.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 354.1490 309.2940 354.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 355.0490 309.2940 355.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 359.5490 309.2940 359.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 357.7500 309.2940 358.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 356.8500 309.2940 357.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 358.6500 309.2940 358.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 355.9500 309.2940 356.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 360.4490 309.2940 360.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 361.3490 309.2940 361.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 364.9500 309.2940 365.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 364.0490 309.2940 364.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 363.1500 309.2940 363.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 362.2490 309.2940 362.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 365.8490 309.2940 366.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 368.5490 309.2940 368.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 367.6500 309.2940 367.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 369.4500 309.2940 369.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 366.7490 309.2940 367.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 373.0500 309.2940 373.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 373.9500 309.2940 374.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 370.3490 309.2940 370.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 374.8500 309.2940 375.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 371.2490 309.2940 371.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 372.1500 309.2940 372.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 375.7490 309.2940 376.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 377.5490 309.2940 377.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 379.3500 309.2940 379.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 376.6490 309.2940 376.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 378.4490 309.2940 378.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 382.0490 309.2940 382.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 381.1500 309.2940 381.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 380.2490 309.2940 380.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 383.8500 309.2940 384.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 382.9490 309.2940 383.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 389.2500 309.2940 389.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 384.7490 309.2940 385.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 385.6500 309.2940 385.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 386.5490 309.2940 386.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 387.4490 309.2940 387.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 388.3500 309.2940 388.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 391.9490 309.2940 392.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 393.7490 309.2940 394.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 390.1500 309.2940 390.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 391.0500 309.2940 391.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 392.8490 309.2940 393.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 398.2490 309.2940 398.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 397.3500 309.2940 397.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 396.4490 309.2940 396.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 395.5500 309.2940 395.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 394.6490 309.2940 394.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 400.9490 309.2940 401.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 400.0500 309.2940 400.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 401.8500 309.2940 402.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 402.7490 309.2940 403.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 399.1490 309.2940 399.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 403.6490 309.2940 403.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 408.1490 309.2940 408.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 405.4500 309.2940 405.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 406.3500 309.2940 406.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 407.2500 309.2940 407.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 404.5500 309.2940 404.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 409.9490 309.2940 410.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 412.6490 309.2940 412.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 411.7500 309.2940 412.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 409.0490 309.2940 409.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 410.8490 309.2940 411.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 414.4490 309.2940 414.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 413.5500 309.2940 413.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 417.1490 309.2940 417.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 416.2500 309.2940 416.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 418.0500 309.2940 418.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 415.3490 309.2940 415.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 421.6500 309.2940 421.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 422.5500 309.2940 422.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 418.9490 309.2940 419.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 419.8490 309.2940 420.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 420.7500 309.2940 421.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 424.3490 309.2940 424.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 426.1490 309.2940 426.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 423.4500 309.2940 423.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 425.2490 309.2940 425.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 427.0490 309.2940 427.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 429.7500 309.2940 430.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 428.8490 309.2940 429.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 430.6490 309.2940 430.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 432.4500 309.2940 432.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 427.9500 309.2940 428.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 431.5490 309.2940 431.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 433.3490 309.2940 433.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 434.2500 309.2940 434.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 435.1490 309.2940 435.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 436.0490 309.2940 436.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 436.9500 309.2940 437.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 440.5490 309.2940 440.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 437.8500 309.2940 438.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 438.7500 309.2940 439.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 439.6500 309.2940 439.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 441.4490 309.2940 441.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 442.3490 309.2940 442.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 445.9500 309.2940 446.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 445.0490 309.2940 445.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 446.8490 309.2940 447.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 444.1500 309.2940 444.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 443.2490 309.2940 443.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 449.5490 309.2940 449.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 448.6500 309.2940 448.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 450.4500 309.2940 450.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 451.3490 309.2940 451.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 447.7490 309.2940 448.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 456.7490 309.2940 457.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 454.0500 309.2940 454.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 454.9500 309.2940 455.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 455.8500 309.2940 456.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 452.2490 309.2940 452.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 453.1500 309.2940 453.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 458.5490 309.2940 458.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 461.2490 309.2940 461.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 460.3500 309.2940 460.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 457.6490 309.2940 457.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 459.4490 309.2940 459.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 462.1500 309.2940 462.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 465.7490 309.2940 466.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 463.0490 309.2940 463.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 464.8500 309.2940 465.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 463.9490 309.2940 464.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 470.2500 309.2940 470.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 471.1500 309.2940 471.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 466.6500 309.2940 466.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 467.5490 309.2940 467.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 468.4490 309.2940 468.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 469.3500 309.2940 469.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 472.9490 309.2940 473.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 474.7490 309.2940 475.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 472.0500 309.2940 472.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 473.8490 309.2940 474.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 475.6490 309.2940 475.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 478.3500 309.2940 478.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 477.4490 309.2940 477.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 479.2490 309.2940 479.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 476.5500 309.2940 476.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 480.1490 309.2940 480.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 481.9490 309.2940 482.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 481.0500 309.2940 481.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 482.8500 309.2940 483.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 483.7490 309.2940 484.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 484.6490 309.2940 484.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 485.5500 309.2940 485.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 489.1490 309.2940 489.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 486.4500 309.2940 486.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 487.3500 309.2940 487.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 488.2500 309.2940 488.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 490.0490 309.2940 490.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 490.9490 309.2940 491.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 494.5500 309.2940 494.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 493.6490 309.2940 493.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 492.7500 309.2940 493.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 491.8490 309.2940 492.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 495.4490 309.2940 495.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 497.2500 309.2940 497.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 499.0500 309.2940 499.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 498.1490 309.2940 498.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 499.9490 309.2940 500.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 496.3490 309.2940 496.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 502.6500 309.2940 502.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 503.5500 309.2940 503.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 504.4500 309.2940 504.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 500.8490 309.2940 501.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 501.7500 309.2940 502.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 505.3490 309.2940 505.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 507.1490 309.2940 507.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 508.9500 309.2940 509.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 506.2490 309.2940 506.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 508.0490 309.2940 508.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 510.7500 309.2940 511.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 509.8490 309.2940 510.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 511.6490 309.2940 511.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 513.4500 309.2940 513.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 514.3490 309.2940 514.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 512.5490 309.2940 512.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 518.8500 309.2940 519.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 515.2500 309.2940 515.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 516.1490 309.2940 516.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 517.0490 309.2940 517.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 517.9500 309.2940 518.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 521.5490 309.2940 521.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 523.3490 309.2940 523.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 519.7500 309.2940 520.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 520.6500 309.2940 520.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 522.4490 309.2940 522.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 526.9500 309.2940 527.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 526.0490 309.2940 526.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 527.8490 309.2940 528.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 525.1500 309.2940 525.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 528.7490 309.2940 529.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 524.2490 309.2940 524.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 529.6500 309.2940 529.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 531.4500 309.2940 531.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 530.5490 309.2940 530.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 532.3490 309.2940 532.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 533.2490 309.2940 533.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 537.7490 309.2940 538.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 535.0500 309.2940 535.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 535.9500 309.2940 536.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 536.8500 309.2940 537.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 534.1500 309.2940 534.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 539.5490 309.2940 539.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 543.1500 309.2940 543.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 542.2490 309.2940 542.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 541.3500 309.2940 541.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 538.6490 309.2940 538.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 540.4490 309.2940 540.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 544.0490 309.2940 544.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 545.8500 309.2940 546.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 547.6500 309.2940 547.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 546.7490 309.2940 547.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 544.9490 309.2940 545.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 551.2500 309.2940 551.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 552.1500 309.2940 552.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 548.5490 309.2940 548.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 553.0500 309.2940 553.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 549.4490 309.2940 549.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 550.3500 309.2940 550.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 553.9490 309.2940 554.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 555.7490 309.2940 556.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 557.5500 309.2940 557.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 554.8490 309.2940 555.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 556.6490 309.2940 556.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 559.3500 309.2940 559.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 558.4490 309.2940 558.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 560.2490 309.2940 560.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 562.0500 309.2940 562.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 561.1490 309.2940 561.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 567.4500 309.2940 567.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 563.8500 309.2940 564.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 562.9490 309.2940 563.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 564.7490 309.2940 565.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 565.6490 309.2940 565.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 566.5500 309.2940 566.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 570.1490 309.2940 570.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 571.9490 309.2940 572.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 568.3500 309.2940 568.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 569.2500 309.2940 569.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 571.0490 309.2940 571.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 575.5500 309.2940 575.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 574.6490 309.2940 574.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 576.4490 309.2940 576.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 573.7500 309.2940 574.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 572.8490 309.2940 573.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 580.0500 309.2940 580.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 579.1490 309.2940 579.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 580.9490 309.2940 581.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 578.2500 309.2940 578.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 577.3490 309.2940 577.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 581.8490 309.2940 582.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 586.3490 309.2940 586.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 583.6500 309.2940 583.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 584.5500 309.2940 584.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 585.4500 309.2940 585.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 582.7500 309.2940 583.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 588.1490 309.2940 588.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 590.8490 309.2940 591.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 589.9500 309.2940 590.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 587.2490 309.2940 587.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 589.0490 309.2940 589.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 591.7500 309.2940 592.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 592.6490 309.2940 592.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 596.2500 309.2940 596.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 595.3490 309.2940 595.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 594.4500 309.2940 594.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 593.5490 309.2940 593.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 599.8500 309.2940 600.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 600.7500 309.2940 601.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 597.1490 309.2940 597.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 598.0490 309.2940 598.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 598.9500 309.2940 599.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 602.5490 309.2940 602.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 604.3490 309.2940 604.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 601.6500 309.2940 601.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 603.4490 309.2940 603.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 605.2490 309.2940 605.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 607.9500 309.2940 608.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 607.0490 309.2940 607.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 608.8490 309.2940 609.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 606.1500 309.2940 606.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 610.6500 309.2940 610.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 609.7490 309.2940 610.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 612.4500 309.2940 612.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 611.5490 309.2940 611.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 613.3490 309.2940 613.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 614.2490 309.2940 614.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 615.1500 309.2940 615.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 618.7490 309.2940 619.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 616.0500 309.2940 616.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 616.9500 309.2940 617.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 617.8500 309.2940 618.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 619.6490 309.2940 619.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 620.5490 309.2940 620.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 624.1500 309.2940 624.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 623.2490 309.2940 623.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 625.0490 309.2940 625.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 622.3500 309.2940 622.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 621.4490 309.2940 621.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 628.6500 309.2940 628.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 627.7490 309.2940 628.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 629.5490 309.2940 629.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 626.8500 309.2940 627.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 625.9490 309.2940 626.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 634.9490 309.2940 635.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 632.2500 309.2940 632.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 633.1500 309.2940 633.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 634.0500 309.2940 634.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 630.4490 309.2940 630.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 631.3500 309.2940 631.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 636.7490 309.2940 637.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 639.4490 309.2940 639.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 638.5500 309.2940 638.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 635.8490 309.2940 636.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 637.6490 309.2940 637.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 640.3500 309.2940 640.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 641.2490 309.2940 641.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 643.9490 309.2940 644.2480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 643.0500 309.2940 643.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 642.1490 309.2940 642.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 648.4500 309.2940 648.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 649.3500 309.2940 649.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 644.8500 309.2940 645.1510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 645.7490 309.2940 646.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 646.6490 309.2940 646.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 647.5500 309.2940 647.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 651.1490 309.2940 651.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 652.9490 309.2940 653.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 650.2500 309.2940 650.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 652.0490 309.2940 652.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 653.8490 309.2940 654.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 656.5500 309.2940 656.8510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 655.6490 309.2940 655.9480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 657.4490 309.2940 657.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 654.7500 309.2940 655.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 658.3490 309.2940 658.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 661.0500 309.2940 661.3510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 660.1490 309.2940 660.4480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 659.2500 309.2940 659.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 661.9490 309.2940 662.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 662.8490 309.2940 663.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 663.7500 309.2940 664.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 667.3490 309.2940 667.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 664.6500 309.2940 664.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 665.5500 309.2940 665.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 666.4500 309.2940 666.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 668.2490 309.2940 668.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 669.1490 309.2940 669.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 672.7500 309.2940 673.0510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 671.8490 309.2940 672.1480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 670.9500 309.2940 671.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 670.0490 309.2940 670.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 673.6490 309.2940 673.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 677.2500 309.2940 677.5510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 676.3490 309.2940 676.6480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 675.4500 309.2940 675.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 674.5490 309.2940 674.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 678.1490 309.2940 678.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 680.8500 309.2940 681.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 681.7500 309.2940 682.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 682.6500 309.2940 682.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 679.0490 309.2940 679.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 679.9500 309.2940 680.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 683.5490 309.2940 683.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 685.3490 309.2940 685.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 687.1500 309.2940 687.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 684.4490 309.2940 684.7500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 686.2490 309.2940 686.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 688.9500 309.2940 689.2510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 688.0490 309.2940 688.3480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 689.8490 309.2940 690.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 692.5490 309.2940 692.8480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 691.6500 309.2940 691.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 690.7490 309.2940 691.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 697.0500 309.2940 697.3500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 693.4500 309.2940 693.7510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 694.3490 309.2940 694.6490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 695.2490 309.2940 695.5490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 696.1500 309.2940 696.4500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 699.7490 309.2940 700.0500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 701.5490 309.2940 701.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 697.9500 309.2940 698.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 698.8500 309.2940 699.1490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 700.6490 309.2940 700.9500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 705.1500 309.2940 705.4510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 704.2490 309.2940 704.5480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 706.0490 309.2940 706.3490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 703.3500 309.2940 703.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 706.9490 309.2940 707.2490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 702.4490 309.2940 702.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 709.6500 309.2940 709.9510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 708.7490 309.2940 709.0480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 707.8500 309.2940 708.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 710.5490 309.2940 710.8490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 711.4490 309.2940 711.7490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 715.9490 309.2940 716.2500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 713.2500 309.2940 713.5500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 714.1500 309.2940 714.4490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 712.3500 309.2940 712.6500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 718.6490 309.2940 718.9490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 716.8490 309.2940 717.1500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 719.5500 309.2940 719.8500 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 720.4490 309.2940 720.7480 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 721.3500 309.2940 721.6510 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 717.7490 309.2940 718.0490 309.5940 ;
    END
    PORT
      LAYER M5 ;
        RECT 715.0500 309.2940 715.3490 309.5940 ;
    END
  END VSS

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 587.6940 0.0000 587.8940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 587.6940 0.0000 587.8940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 587.6940 0.0000 587.8940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 587.6940 0.0000 587.8940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 587.6940 0.0000 587.8940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[44]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 586.3260 0.0000 586.5260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 586.3260 0.0000 586.5260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 586.3260 0.0000 586.5260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 586.3260 0.0000 586.5260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 586.3260 0.0000 586.5260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[43]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 585.6410 0.0000 585.8410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 585.6410 0.0000 585.8410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 585.6410 0.0000 585.8410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 585.6410 0.0000 585.8410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 585.6410 0.0000 585.8410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 589.7450 0.0000 589.9450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 589.7450 0.0000 589.9450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 589.7450 0.0000 589.9450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 589.7450 0.0000 589.9450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 589.7450 0.0000 589.9450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[46]

  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 590.4300 0.0000 590.6300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 590.4300 0.0000 590.6300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 590.4300 0.0000 590.6300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 590.4300 0.0000 590.6300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 590.4300 0.0000 590.6300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[46]

  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 591.1130 0.0010 591.3130 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 591.1130 0.0010 591.3130 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 591.1130 0.0000 591.3130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 591.1130 0.0000 591.3130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 591.1130 0.0000 591.3130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[47]

  PIN I[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 593.8490 0.0000 594.0490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 593.8490 0.0000 594.0490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 593.8490 0.0000 594.0490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 593.8490 0.0000 594.0490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 593.8490 0.0000 594.0490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[49]

  PIN O[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 594.5340 0.0000 594.7340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 594.5340 0.0000 594.7340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 594.5340 0.0000 594.7340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 594.5340 0.0000 594.7340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 594.5340 0.0000 594.7340 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[49]

  PIN I[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 595.2170 0.0000 595.4170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 595.2170 0.0000 595.4170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 595.2170 0.0000 595.4170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 595.2170 0.0000 595.4170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 595.2170 0.0000 595.4170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[50]

  PIN O[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 595.9020 0.0000 596.1020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 595.9020 0.0000 596.1020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 595.9020 0.0000 596.1020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 595.9020 0.0000 596.1020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 595.9020 0.0000 596.1020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[50]

  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 591.7980 0.0000 591.9980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 591.7980 0.0000 591.9980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 591.7980 0.0000 591.9980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 591.7980 0.0000 591.9980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 591.7980 0.0000 591.9980 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[47]

  PIN O[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 593.1660 0.0000 593.3660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 593.1660 0.0000 593.3660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 593.1660 0.0000 593.3660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 593.1660 0.0000 593.3660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 593.1660 0.0000 593.3660 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[48]

  PIN I[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 592.4810 0.0000 592.6810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 592.4810 0.0000 592.6810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 592.4810 0.0000 592.6810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 592.4810 0.0000 592.6810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 592.4810 0.0000 592.6810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[48]

  PIN I[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 596.5850 0.0000 596.7850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 596.5850 0.0000 596.7850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 596.5850 0.0000 596.7850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 596.5850 0.0000 596.7850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 596.5850 0.0000 596.7850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[51]

  PIN O[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 597.2700 0.0000 597.4700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 597.2700 0.0000 597.4700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 597.2700 0.0000 597.4700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 597.2700 0.0000 597.4700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 597.2700 0.0000 597.4700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[51]

  PIN O[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 600.0060 0.0000 600.2060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 600.0060 0.0000 600.2060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 600.0060 0.0000 600.2060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 600.0060 0.0000 600.2060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 600.0060 0.0000 600.2060 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[53]

  PIN O[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 601.3740 0.0000 601.5740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 601.3740 0.0000 601.5740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 601.3740 0.0000 601.5740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 601.3740 0.0000 601.5740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 601.3740 0.0000 601.5740 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[54]

  PIN I[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 600.6890 0.0000 600.8890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 600.6890 0.0000 600.8890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 600.6890 0.0000 600.8890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 600.6890 0.0000 600.8890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 600.6890 0.0000 600.8890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[54]

  PIN I[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 602.0570 0.0000 602.2570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 602.0570 0.0000 602.2570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 602.0570 0.0000 602.2570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 602.0570 0.0000 602.2570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 602.0570 0.0000 602.2570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[55]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 575.3820 0.0000 575.5820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 575.3820 0.0000 575.5820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 575.3820 0.0000 575.5820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 575.3820 0.0000 575.5820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 575.3820 0.0000 575.5820 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[35]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 576.0650 0.0000 576.2650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 576.0650 0.0000 576.2650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 576.0650 0.0000 576.2650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 576.0650 0.0000 576.2650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 576.0650 0.0000 576.2650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 576.7500 0.0000 576.9500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 576.7500 0.0000 576.9500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 576.7500 0.0000 576.9500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 576.7500 0.0000 576.9500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 576.7500 0.0000 576.9500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[36]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 574.6970 0.0000 574.8970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 574.6970 0.0000 574.8970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 574.6970 0.0000 574.8970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 574.6970 0.0000 574.8970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 574.6970 0.0000 574.8970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 573.3290 0.0000 573.5290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 573.3290 0.0000 573.5290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 573.3290 0.0000 573.5290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 573.3290 0.0000 573.5290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 573.3290 0.0000 573.5290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 574.0140 0.0000 574.2140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 574.0140 0.0000 574.2140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 574.0140 0.0000 574.2140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 574.0140 0.0000 574.2140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 574.0140 0.0000 574.2140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[34]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 578.8010 0.0000 579.0010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 578.8010 0.0000 579.0010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 578.8010 0.0000 579.0010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 578.8010 0.0000 579.0010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 578.8010 0.0000 579.0010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 582.2220 0.0000 582.4220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 582.2220 0.0000 582.4220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 582.2220 0.0000 582.4220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 582.2220 0.0000 582.4220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 582.2220 0.0000 582.4220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[40]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 580.1690 0.0000 580.3690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 580.1690 0.0000 580.3690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 580.1690 0.0000 580.3690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 580.1690 0.0000 580.3690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 580.1690 0.0000 580.3690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[39]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 581.5370 0.0000 581.7370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 581.5370 0.0000 581.7370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 581.5370 0.0000 581.7370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 581.5370 0.0000 581.7370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 581.5370 0.0000 581.7370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[40]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 580.8540 0.0000 581.0540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 580.8540 0.0000 581.0540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 580.8540 0.0000 581.0540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 580.8540 0.0000 581.0540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 580.8540 0.0000 581.0540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[39]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 579.4860 0.0000 579.6860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 579.4860 0.0000 579.6860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 579.4860 0.0000 579.6860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 579.4860 0.0000 579.6860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 579.4860 0.0000 579.6860 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[38]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 584.9580 0.0000 585.1580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 584.9580 0.0000 585.1580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 584.9580 0.0000 585.1580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 584.9580 0.0000 585.1580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 584.9580 0.0000 585.1580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[42]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 584.2730 0.0000 584.4730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 584.2730 0.0000 584.4730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 584.2730 0.0000 584.4730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 584.2730 0.0000 584.4730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 584.2730 0.0000 584.4730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[42]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 583.5900 0.0000 583.7900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 583.5900 0.0000 583.7900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 583.5900 0.0000 583.7900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 583.5900 0.0000 583.7900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 583.5900 0.0000 583.7900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[41]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 582.9050 0.0000 583.1050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 582.9050 0.0000 583.1050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 582.9050 0.0000 583.1050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 582.9050 0.0000 583.1050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 582.9050 0.0000 583.1050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[41]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 588.3770 0.0000 588.5770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 588.3770 0.0000 588.5770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 588.3770 0.0000 588.5770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 588.3770 0.0000 588.5770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 588.3770 0.0000 588.5770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 589.0620 0.0000 589.2620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 589.0620 0.0000 589.2620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 589.0620 0.0000 589.2620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 589.0620 0.0000 589.2620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 589.0620 0.0000 589.2620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[45]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 563.0700 0.0000 563.2700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 563.0700 0.0000 563.2700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 563.0700 0.0000 563.2700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 563.0700 0.0000 563.2700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 563.0700 0.0000 563.2700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[26]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 561.7020 0.0000 561.9020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 561.7020 0.0000 561.9020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 561.7020 0.0000 561.9020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 561.7020 0.0000 561.9020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 561.7020 0.0000 561.9020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[25]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 561.0170 0.0000 561.2170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 561.0170 0.0000 561.2170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 561.0170 0.0000 561.2170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 561.0170 0.0000 561.2170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 561.0170 0.0000 561.2170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 566.4890 0.0000 566.6890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 566.4890 0.0000 566.6890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 566.4890 0.0000 566.6890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 566.4890 0.0000 566.6890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 566.4890 0.0000 566.6890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 565.8060 0.0000 566.0060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 565.8060 0.0000 566.0060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 565.8060 0.0000 566.0060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 565.8060 0.0000 566.0060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 565.8060 0.0000 566.0060 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[28]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 565.1210 0.0000 565.3210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 565.1210 0.0000 565.3210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 565.1210 0.0000 565.3210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 565.1210 0.0000 565.3210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 565.1210 0.0000 565.3210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 563.7530 0.0000 563.9530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 563.7530 0.0000 563.9530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 563.7530 0.0000 563.9530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 563.7530 0.0000 563.9530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 563.7530 0.0000 563.9530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 564.4380 0.0000 564.6380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 564.4380 0.0000 564.6380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 564.4380 0.0000 564.6380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 564.4380 0.0000 564.6380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 564.4380 0.0000 564.6380 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[27]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 569.9100 0.0000 570.1100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 569.9100 0.0000 570.1100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 569.9100 0.0000 570.1100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 569.9100 0.0000 570.1100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 569.9100 0.0000 570.1100 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[31]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 569.2250 0.0000 569.4250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 569.2250 0.0000 569.4250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 569.2250 0.0000 569.4250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 569.2250 0.0000 569.4250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 569.2250 0.0000 569.4250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 568.5420 0.0000 568.7420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 568.5420 0.0000 568.7420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 568.5420 0.0000 568.7420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 568.5420 0.0000 568.7420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 568.5420 0.0000 568.7420 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[30]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 567.8570 0.0000 568.0570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 567.8570 0.0000 568.0570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 567.8570 0.0000 568.0570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 567.8570 0.0000 568.0570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 567.8570 0.0000 568.0570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 567.1740 0.0000 567.3740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 567.1740 0.0000 567.3740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 567.1740 0.0000 567.3740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 567.1740 0.0000 567.3740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 567.1740 0.0000 567.3740 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[29]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 572.6460 0.0000 572.8460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 572.6460 0.0000 572.8460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 572.6460 0.0000 572.8460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 572.6460 0.0000 572.8460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 572.6460 0.0000 572.8460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[33]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 571.9610 0.0000 572.1610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 571.9610 0.0000 572.1610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 571.9610 0.0000 572.1610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 571.9610 0.0000 572.1610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 571.9610 0.0000 572.1610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 570.5930 0.0000 570.7930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 570.5930 0.0000 570.7930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 570.5930 0.0000 570.7930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 570.5930 0.0000 570.7930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 570.5930 0.0000 570.7930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 571.2780 0.0000 571.4780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 571.2780 0.0000 571.4780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 571.2780 0.0000 571.4780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 571.2780 0.0000 571.4780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 571.2780 0.0000 571.4780 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[32]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 577.4330 0.0000 577.6330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 577.4330 0.0000 577.6330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 577.4330 0.0000 577.6330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 577.4330 0.0000 577.6330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 577.4330 0.0000 577.6330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[37]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 578.1180 0.0000 578.3180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 578.1180 0.0000 578.3180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 578.1180 0.0000 578.3180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 578.1180 0.0000 578.3180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 578.1180 0.0000 578.3180 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[37]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 548.7050 0.0000 548.9050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 548.7050 0.0000 548.9050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 548.7050 0.0000 548.9050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 548.7050 0.0000 548.9050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 548.7050 0.0000 548.9050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 549.3900 0.0000 549.5900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 549.3900 0.0000 549.5900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 549.3900 0.0000 549.5900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 549.3900 0.0000 549.5900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 549.3900 0.0000 549.5900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[16]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 550.0730 0.0000 550.2730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 550.0730 0.0000 550.2730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 550.0730 0.0000 550.2730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 550.0730 0.0000 550.2730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 550.0730 0.0000 550.2730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 553.4940 0.0000 553.6940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 553.4940 0.0000 553.6940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 553.4940 0.0000 553.6940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 553.4940 0.0000 553.6940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 553.4940 0.0000 553.6940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[19]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 554.1770 0.0000 554.3770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 554.1770 0.0000 554.3770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 554.1770 0.0000 554.3770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 554.1770 0.0000 554.3770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 554.1770 0.0000 554.3770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 552.8090 0.0000 553.0090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 552.8090 0.0000 553.0090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 552.8090 0.0000 553.0090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 552.8090 0.0000 553.0090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 552.8090 0.0000 553.0090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 552.1260 0.0000 552.3260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 552.1260 0.0000 552.3260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 552.1260 0.0000 552.3260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 552.1260 0.0000 552.3260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 552.1260 0.0000 552.3260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[18]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 551.4410 0.0000 551.6410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 551.4410 0.0000 551.6410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 551.4410 0.0000 551.6410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 551.4410 0.0000 551.6410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 551.4410 0.0000 551.6410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 557.5980 0.0000 557.7980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 557.5980 0.0000 557.7980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 557.5980 0.0000 557.7980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 557.5980 0.0000 557.7980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 557.5980 0.0000 557.7980 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[22]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 556.9130 0.0000 557.1130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 556.9130 0.0000 557.1130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 556.9130 0.0000 557.1130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 556.9130 0.0000 557.1130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 556.9130 0.0000 557.1130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 555.5450 0.0000 555.7450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 555.5450 0.0000 555.7450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 555.5450 0.0000 555.7450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 555.5450 0.0000 555.7450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 555.5450 0.0000 555.7450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 556.2300 0.0000 556.4300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 556.2300 0.0000 556.4300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 556.2300 0.0000 556.4300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 556.2300 0.0000 556.4300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 556.2300 0.0000 556.4300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[21]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 554.8620 0.0000 555.0620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 554.8620 0.0000 555.0620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 554.8620 0.0000 555.0620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 554.8620 0.0000 555.0620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 554.8620 0.0000 555.0620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[20]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 558.9660 0.0000 559.1660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 558.9660 0.0000 559.1660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 558.9660 0.0000 559.1660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 558.9660 0.0000 559.1660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 558.9660 0.0000 559.1660 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[23]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 559.6490 0.0000 559.8490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 559.6490 0.0000 559.8490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 559.6490 0.0000 559.8490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 559.6490 0.0000 559.8490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 559.6490 0.0000 559.8490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 560.3340 0.0000 560.5340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 560.3340 0.0000 560.5340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 560.3340 0.0000 560.5340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 560.3340 0.0000 560.5340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 560.3340 0.0000 560.5340 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[24]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 558.2810 0.0000 558.4810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 558.2810 0.0000 558.4810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 558.2810 0.0000 558.4810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 558.2810 0.0000 558.4810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 558.2810 0.0000 558.4810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 562.3850 0.0000 562.5850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 562.3850 0.0000 562.5850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 562.3850 0.0000 562.5850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 562.3850 0.0000 562.5850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 562.3850 0.0000 562.5850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 536.3930 0.0000 536.5930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 536.3930 0.0000 536.5930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 536.3930 0.0000 536.5930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 536.3930 0.0000 536.5930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 536.3930 0.0000 536.5930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 541.8650 0.0000 542.0650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 541.8650 0.0000 542.0650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 541.8650 0.0000 542.0650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 541.8650 0.0000 542.0650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 541.8650 0.0000 542.0650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 540.4970 0.0000 540.6970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 540.4970 0.0000 540.6970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 540.4970 0.0000 540.6970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 540.4970 0.0000 540.6970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 540.4970 0.0000 540.6970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 541.1820 0.0000 541.3820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 541.1820 0.0000 541.3820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 541.1820 0.0000 541.3820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 541.1820 0.0000 541.3820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 541.1820 0.0000 541.3820 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[10]

  PIN O[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 660.1980 0.0000 660.3980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 660.1980 0.0000 660.3980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 660.1980 0.0000 660.3980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 660.1980 0.0000 660.3980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 660.1980 0.0000 660.3980 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[97]

  PIN O[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 665.6700 0.0000 665.8700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 665.6700 0.0000 665.8700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 665.6700 0.0000 665.8700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 665.6700 0.0000 665.8700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 665.6700 0.0000 665.8700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[101]

  PIN I[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 664.9850 0.0000 665.1850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 664.9850 0.0000 665.1850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 664.9850 0.0000 665.1850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 664.9850 0.0000 665.1850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 664.9850 0.0000 665.1850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[101]

  PIN O[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.6780 0.0000 639.8780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 639.6780 0.0000 639.8780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 639.6780 0.0000 639.8780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 639.6780 0.0000 639.8780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 639.6780 0.0000 639.8780 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[82]

  PIN I[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 638.9930 0.0000 639.1930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 638.9930 0.0000 639.1930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 638.9930 0.0000 639.1930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 638.9930 0.0000 639.1930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 638.9930 0.0000 639.1930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[82]

  PIN O[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 641.0460 0.0000 641.2460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 641.0460 0.0000 641.2460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 641.0460 0.0000 641.2460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 641.0460 0.0000 641.2460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 641.0460 0.0000 641.2460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[83]

  PIN I[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 640.3610 0.0000 640.5610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 640.3610 0.0000 640.5610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 640.3610 0.0000 640.5610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 640.3610 0.0000 640.5610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 640.3610 0.0000 640.5610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[83]

  PIN I[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 641.7290 0.0000 641.9290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 641.7290 0.0000 641.9290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 641.7290 0.0000 641.9290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 641.7290 0.0000 641.9290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 641.7290 0.0000 641.9290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[84]

  PIN O[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 643.7820 0.0000 643.9820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 643.7820 0.0000 643.9820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 643.7820 0.0000 643.9820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 643.7820 0.0000 643.9820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 643.7820 0.0000 643.9820 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[85]

  PIN I[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 644.4650 0.0000 644.6650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 644.4650 0.0000 644.6650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 644.4650 0.0000 644.6650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 644.4650 0.0000 644.6650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 644.4650 0.0000 644.6650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[86]

  PIN I[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 643.0970 0.0000 643.2970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 643.0970 0.0000 643.2970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 643.0970 0.0000 643.2970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 643.0970 0.0000 643.2970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 643.0970 0.0000 643.2970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[85]

  PIN O[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 645.1500 0.0000 645.3500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 645.1500 0.0000 645.3500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 645.1500 0.0000 645.3500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 645.1500 0.0000 645.3500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 645.1500 0.0000 645.3500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[86]

  PIN O[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 642.4140 0.0000 642.6140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 642.4140 0.0000 642.6140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 642.4140 0.0000 642.6140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 642.4140 0.0000 642.6140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 642.4140 0.0000 642.6140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[84]

  PIN I[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 645.8330 0.0000 646.0330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 645.8330 0.0000 646.0330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 645.8330 0.0000 646.0330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 645.8330 0.0000 646.0330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 645.8330 0.0000 646.0330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[87]

  PIN O[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 646.5180 0.0000 646.7180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 646.5180 0.0000 646.7180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 646.5180 0.0000 646.7180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 646.5180 0.0000 646.7180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 646.5180 0.0000 646.7180 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[87]

  PIN I[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 647.2010 0.0000 647.4010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 647.2010 0.0000 647.4010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 647.2010 0.0000 647.4010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 647.2010 0.0000 647.4010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 647.2010 0.0000 647.4010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[88]

  PIN O[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 649.2540 0.0000 649.4540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 649.2540 0.0000 649.4540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 649.2540 0.0000 649.4540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 649.2540 0.0000 649.4540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 649.2540 0.0000 649.4540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[89]

  PIN O[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 650.6220 0.0000 650.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 650.6220 0.0000 650.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 650.6220 0.0000 650.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 650.6220 0.0000 650.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 650.6220 0.0000 650.8220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[90]

  PIN I[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 649.9370 0.0000 650.1370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 649.9370 0.0000 650.1370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 649.9370 0.0000 650.1370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 649.9370 0.0000 650.1370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 649.9370 0.0000 650.1370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[90]

  PIN I[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 648.5690 0.0000 648.7690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 648.5690 0.0000 648.7690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 648.5690 0.0000 648.7690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 648.5690 0.0000 648.7690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 648.5690 0.0000 648.7690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[89]

  PIN O[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 647.8860 0.0000 648.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 647.8860 0.0000 648.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 647.8860 0.0000 648.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 647.8860 0.0000 648.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 647.8860 0.0000 648.0860 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[88]

  PIN O[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 623.2620 0.0000 623.4620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 623.2620 0.0000 623.4620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 623.2620 0.0000 623.4620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 623.2620 0.0000 623.4620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 623.2620 0.0000 623.4620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[70]

  PIN I[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 623.9450 0.0000 624.1450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 623.9450 0.0000 624.1450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 623.9450 0.0000 624.1450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 623.9450 0.0000 624.1450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 623.9450 0.0000 624.1450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[71]

  PIN O[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 627.3660 0.0000 627.5660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 627.3660 0.0000 627.5660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 627.3660 0.0000 627.5660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 627.3660 0.0000 627.5660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 627.3660 0.0000 627.5660 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[73]

  PIN I[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 628.0490 0.0000 628.2490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 628.0490 0.0000 628.2490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 628.0490 0.0000 628.2490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 628.0490 0.0000 628.2490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 628.0490 0.0000 628.2490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[74]

  PIN O[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 628.7340 0.0000 628.9340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 628.7340 0.0000 628.9340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 628.7340 0.0000 628.9340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 628.7340 0.0000 628.9340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 628.7340 0.0000 628.9340 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[74]

  PIN O[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 630.1020 0.0000 630.3020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 630.1020 0.0000 630.3020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 630.1020 0.0000 630.3020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 630.1020 0.0000 630.3020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 630.1020 0.0000 630.3020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[75]

  PIN I[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 629.4170 0.0000 629.6170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 629.4170 0.0000 629.6170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 629.4170 0.0000 629.6170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 629.4170 0.0000 629.6170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 629.4170 0.0000 629.6170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[75]

  PIN I[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 630.7850 0.0000 630.9850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 630.7850 0.0000 630.9850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 630.7850 0.0000 630.9850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 630.7850 0.0000 630.9850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 630.7850 0.0000 630.9850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[76]

  PIN O[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 631.4700 0.0000 631.6700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 631.4700 0.0000 631.6700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 631.4700 0.0000 631.6700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 631.4700 0.0000 631.6700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 631.4700 0.0000 631.6700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[76]

  PIN I[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 632.1530 0.0000 632.3530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 632.1530 0.0000 632.3530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 632.1530 0.0000 632.3530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 632.1530 0.0000 632.3530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 632.1530 0.0000 632.3530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[77]

  PIN O[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 632.8380 0.0000 633.0380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 632.8380 0.0000 633.0380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 632.8380 0.0000 633.0380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 632.8380 0.0000 633.0380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 632.8380 0.0000 633.0380 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[77]

  PIN O[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 634.2060 0.0000 634.4060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 634.2060 0.0000 634.4060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 634.2060 0.0000 634.4060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 634.2060 0.0000 634.4060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 634.2060 0.0000 634.4060 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[78]

  PIN I[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 633.5210 0.0000 633.7210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 633.5210 0.0000 633.7210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 633.5210 0.0000 633.7210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 633.5210 0.0000 633.7210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 633.5210 0.0000 633.7210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[78]

  PIN I[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 634.8890 0.0000 635.0890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 634.8890 0.0000 635.0890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 634.8890 0.0000 635.0890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 634.8890 0.0000 635.0890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 634.8890 0.0000 635.0890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[79]

  PIN O[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 636.9420 0.0000 637.1420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 636.9420 0.0000 637.1420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 636.9420 0.0000 637.1420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 636.9420 0.0000 637.1420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 636.9420 0.0000 637.1420 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[80]

  PIN I[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 637.6250 0.0000 637.8250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 637.6250 0.0000 637.8250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 637.6250 0.0000 637.8250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 637.6250 0.0000 637.8250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 637.6250 0.0000 637.8250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[81]

  PIN O[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 638.3100 0.0000 638.5100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 638.3100 0.0000 638.5100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 638.3100 0.0000 638.5100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 638.3100 0.0000 638.5100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 638.3100 0.0000 638.5100 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[81]

  PIN O[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 635.5740 0.0000 635.7740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 635.5740 0.0000 635.7740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 635.5740 0.0000 635.7740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 635.5740 0.0000 635.7740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 635.5740 0.0000 635.7740 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[79]

  PIN I[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 636.2570 0.0000 636.4570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 636.2570 0.0000 636.4570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 636.2570 0.0000 636.4570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 636.2570 0.0000 636.4570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 636.2570 0.0000 636.4570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[80]

  PIN O[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 610.9500 0.0000 611.1500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 610.9500 0.0000 611.1500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 610.9500 0.0000 611.1500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 610.9500 0.0000 611.1500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 610.9500 0.0000 611.1500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[61]

  PIN I[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 610.2650 0.0000 610.4650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 610.2650 0.0000 610.4650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 610.2650 0.0000 610.4650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 610.2650 0.0000 610.4650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 610.2650 0.0000 610.4650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[61]

  PIN I[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 611.6330 0.0000 611.8330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 611.6330 0.0000 611.8330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 611.6330 0.0000 611.8330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 611.6330 0.0000 611.8330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 611.6330 0.0000 611.8330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[62]

  PIN O[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 615.0540 0.0000 615.2540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 615.0540 0.0000 615.2540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 615.0540 0.0000 615.2540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 615.0540 0.0000 615.2540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 615.0540 0.0000 615.2540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[64]

  PIN I[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 615.7370 0.0000 615.9370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 615.7370 0.0000 615.9370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 615.7370 0.0000 615.9370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 615.7370 0.0000 615.9370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 615.7370 0.0000 615.9370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[65]

  PIN I[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 617.1050 0.0000 617.3050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 617.1050 0.0000 617.3050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 617.1050 0.0000 617.3050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 617.1050 0.0000 617.3050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 617.1050 0.0000 617.3050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[66]

  PIN O[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 616.4220 0.0000 616.6220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 616.4220 0.0000 616.6220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 616.4220 0.0000 616.6220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 616.4220 0.0000 616.6220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 616.4220 0.0000 616.6220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[65]

  PIN O[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 617.7900 0.0000 617.9900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 617.7900 0.0000 617.9900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 617.7900 0.0000 617.9900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 617.7900 0.0000 617.9900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 617.7900 0.0000 617.9900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[66]

  PIN O[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 619.1580 0.0000 619.3580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 619.1580 0.0000 619.3580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 619.1580 0.0000 619.3580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 619.1580 0.0000 619.3580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 619.1580 0.0000 619.3580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[67]

  PIN I[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 618.4730 0.0000 618.6730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 618.4730 0.0000 618.6730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 618.4730 0.0000 618.6730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 618.4730 0.0000 618.6730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 618.4730 0.0000 618.6730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[67]

  PIN I[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 619.8410 0.0000 620.0410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 619.8410 0.0000 620.0410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 619.8410 0.0000 620.0410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 619.8410 0.0000 620.0410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 619.8410 0.0000 620.0410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[68]

  PIN O[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 620.5260 0.0000 620.7260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 620.5260 0.0000 620.7260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 620.5260 0.0000 620.7260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 620.5260 0.0000 620.7260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 620.5260 0.0000 620.7260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[68]

  PIN I[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 621.2090 0.0000 621.4090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 621.2090 0.0000 621.4090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 621.2090 0.0000 621.4090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 621.2090 0.0000 621.4090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 621.2090 0.0000 621.4090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[69]

  PIN I[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 622.5770 0.0000 622.7770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 622.5770 0.0000 622.7770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 622.5770 0.0000 622.7770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 622.5770 0.0000 622.7770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 622.5770 0.0000 622.7770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[70]

  PIN O[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 621.8940 0.0000 622.0940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 621.8940 0.0000 622.0940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 621.8940 0.0000 622.0940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 621.8940 0.0000 622.0940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 621.8940 0.0000 622.0940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[69]

  PIN O[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 624.6300 0.0000 624.8300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 624.6300 0.0000 624.8300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 624.6300 0.0000 624.8300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 624.6300 0.0000 624.8300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 624.6300 0.0000 624.8300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[71]

  PIN O[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 625.9980 0.0000 626.1980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 625.9980 0.0000 626.1980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 625.9980 0.0000 626.1980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 625.9980 0.0000 626.1980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 625.9980 0.0000 626.1980 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[72]

  PIN I[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 625.3130 0.0000 625.5130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 625.3130 0.0000 625.5130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 625.3130 0.0000 625.5130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 625.3130 0.0000 625.5130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 625.3130 0.0000 625.5130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[72]

  PIN I[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 626.6810 0.0000 626.8810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 626.6810 0.0000 626.8810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 626.6810 0.0000 626.8810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 626.6810 0.0000 626.8810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 626.6810 0.0000 626.8810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[73]

  PIN I[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 597.9530 0.0000 598.1530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 597.9530 0.0000 598.1530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 597.9530 0.0000 598.1530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 597.9530 0.0000 598.1530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 597.9530 0.0000 598.1530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[52]

  PIN O[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 598.6380 0.0000 598.8380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 598.6380 0.0000 598.8380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 598.6380 0.0000 598.8380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 598.6380 0.0000 598.8380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 598.6380 0.0000 598.8380 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[52]

  PIN I[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 599.3210 0.0000 599.5210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 599.3210 0.0000 599.5210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 599.3210 0.0000 599.5210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 599.3210 0.0000 599.5210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 599.3210 0.0000 599.5210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[53]

  PIN O[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 602.7420 0.0000 602.9420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 602.7420 0.0000 602.9420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 602.7420 0.0000 602.9420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 602.7420 0.0000 602.9420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 602.7420 0.0000 602.9420 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[55]

  PIN I[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 603.4250 0.0000 603.6250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 603.4250 0.0000 603.6250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 603.4250 0.0000 603.6250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 603.4250 0.0000 603.6250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 603.4250 0.0000 603.6250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[56]

  PIN O[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 604.1100 0.0000 604.3100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 604.1100 0.0000 604.3100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 604.1100 0.0000 604.3100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 604.1100 0.0000 604.3100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 604.1100 0.0000 604.3100 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[56]

  PIN I[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 604.7930 0.0000 604.9930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 604.7930 0.0000 604.9930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 604.7930 0.0000 604.9930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 604.7930 0.0000 604.9930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 604.7930 0.0000 604.9930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[57]

  PIN O[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 605.4780 0.0000 605.6780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 605.4780 0.0000 605.6780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 605.4780 0.0000 605.6780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 605.4780 0.0000 605.6780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 605.4780 0.0000 605.6780 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[57]

  PIN I[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 606.1610 0.0000 606.3610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 606.1610 0.0000 606.3610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 606.1610 0.0000 606.3610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 606.1610 0.0000 606.3610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 606.1610 0.0000 606.3610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[58]

  PIN O[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 606.8460 0.0000 607.0460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 606.8460 0.0000 607.0460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 606.8460 0.0000 607.0460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 606.8460 0.0000 607.0460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 606.8460 0.0000 607.0460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[58]

  PIN O[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 608.2140 0.0000 608.4140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 608.2140 0.0000 608.4140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 608.2140 0.0000 608.4140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 608.2140 0.0000 608.4140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 608.2140 0.0000 608.4140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[59]

  PIN I[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 607.5290 0.0000 607.7290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 607.5290 0.0000 607.7290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 607.5290 0.0000 607.7290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 607.5290 0.0000 607.7290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 607.5290 0.0000 607.7290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[59]

  PIN I[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 608.8970 0.0000 609.0970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 608.8970 0.0000 609.0970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 608.8970 0.0000 609.0970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 608.8970 0.0000 609.0970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 608.8970 0.0000 609.0970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[60]

  PIN O[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 609.5820 0.0000 609.7820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 609.5820 0.0000 609.7820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 609.5820 0.0000 609.7820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 609.5820 0.0000 609.7820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 609.5820 0.0000 609.7820 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[60]

  PIN I[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 613.0010 0.0000 613.2010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 613.0010 0.0000 613.2010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 613.0010 0.0000 613.2010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 613.0010 0.0000 613.2010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 613.0010 0.0000 613.2010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[63]

  PIN O[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 612.3180 0.0000 612.5180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 612.3180 0.0000 612.5180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 612.3180 0.0000 612.5180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 612.3180 0.0000 612.5180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 612.3180 0.0000 612.5180 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[62]

  PIN O[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 613.6860 0.0000 613.8860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 613.6860 0.0000 613.8860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 613.6860 0.0000 613.8860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 613.6860 0.0000 613.8860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 613.6860 0.0000 613.8860 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[63]

  PIN I[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 614.3690 0.0000 614.5690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 614.3690 0.0000 614.5690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 614.3690 0.0000 614.5690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 614.3690 0.0000 614.5690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 614.3690 0.0000 614.5690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[64]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 587.0090 0.0000 587.2090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 587.0090 0.0000 587.2090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 587.0090 0.0000 587.2090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 587.0090 0.0000 587.2090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 587.0090 0.0000 587.2090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 722.9820 245.5700 723.1820 245.7700 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 245.5700 723.1820 245.7700 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 245.5700 723.1820 245.7700 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 245.5700 723.1820 245.7700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 9.8200 723.1820 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 9.8200 723.1820 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 9.8200 723.1820 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 9.8200 723.1820 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 9.8200 723.1820 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 16.8280 723.1820 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 16.8280 723.1820 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 16.8280 723.1820 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 16.8280 723.1820 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 16.8280 723.1820 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9880 288.0560 723.1820 288.2560 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9880 288.0560 723.1820 288.2560 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9880 288.0560 723.1820 288.2560 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9880 288.0560 723.1820 288.2560 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9880 288.0560 723.1820 288.2560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 701.9110 0.0000 702.1110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 701.9110 0.0000 702.1110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 701.9110 0.0000 702.1110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 701.9110 0.0000 702.1110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 701.9110 0.0000 702.1110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 89.4700 723.1820 89.6700 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 89.4700 723.1820 89.6700 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 89.4700 723.1820 89.6700 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 89.4700 723.1820 89.6700 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 89.4700 723.1820 89.6700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 722.9820 89.1090 723.1820 89.3090 ;
    END
    PORT
      LAYER M4 ;
        RECT 722.9820 89.1090 723.1820 89.3090 ;
    END
    PORT
      LAYER M3 ;
        RECT 722.9820 89.1090 723.1820 89.3090 ;
    END
    PORT
      LAYER M2 ;
        RECT 722.9820 89.1090 723.1820 89.3090 ;
    END
    PORT
      LAYER M1 ;
        RECT 722.9820 89.1090 723.1820 89.3090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[8]

  PIN O[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 688.9260 0.0000 689.1260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 688.9260 0.0000 689.1260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 688.9260 0.0000 689.1260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 688.9260 0.0000 689.1260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 688.9260 0.0000 689.1260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[118]

  PIN O[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 687.5580 0.0000 687.7580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 687.5580 0.0000 687.7580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 687.5580 0.0000 687.7580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 687.5580 0.0000 687.7580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 687.5580 0.0000 687.7580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[117]

  PIN I[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 692.3450 0.0000 692.5450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 692.3450 0.0000 692.5450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 692.3450 0.0000 692.5450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 692.3450 0.0000 692.5450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 692.3450 0.0000 692.5450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[121]

  PIN O[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 691.6620 0.0000 691.8620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 691.6620 0.0000 691.8620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 691.6620 0.0000 691.8620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 691.6620 0.0000 691.8620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 691.6620 0.0000 691.8620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[120]

  PIN O[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 693.0300 0.0000 693.2300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 693.0300 0.0000 693.2300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 693.0300 0.0000 693.2300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 693.0300 0.0000 693.2300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 693.0300 0.0000 693.2300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[121]

  PIN I[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 690.9770 0.0000 691.1770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 690.9770 0.0000 691.1770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 690.9770 0.0000 691.1770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 690.9770 0.0000 691.1770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 690.9770 0.0000 691.1770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[120]

  PIN I[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 696.4490 0.0000 696.6490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 696.4490 0.0000 696.6490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 696.4490 0.0000 696.6490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 696.4490 0.0000 696.6490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 696.4490 0.0000 696.6490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[124]

  PIN O[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 695.7660 0.0000 695.9660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 695.7660 0.0000 695.9660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 695.7660 0.0000 695.9660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 695.7660 0.0000 695.9660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 695.7660 0.0000 695.9660 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[123]

  PIN I[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 695.0810 0.0000 695.2810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 695.0810 0.0000 695.2810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 695.0810 0.0000 695.2810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 695.0810 0.0000 695.2810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 695.0810 0.0000 695.2810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[123]

  PIN O[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 694.3980 0.0000 694.5980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 694.3980 0.0000 694.5980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 694.3980 0.0000 694.5980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 694.3980 0.0000 694.5980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 694.3980 0.0000 694.5980 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[122]

  PIN I[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 693.7130 0.0000 693.9130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 693.7130 0.0000 693.9130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 693.7130 0.0000 693.9130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 693.7130 0.0000 693.9130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 693.7130 0.0000 693.9130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[122]

  PIN O[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 698.5020 0.0000 698.7020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 698.5020 0.0000 698.7020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 698.5020 0.0000 698.7020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 698.5020 0.0000 698.7020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 698.5020 0.0000 698.7020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[125]

  PIN I[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 697.8170 0.0000 698.0170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 697.8170 0.0000 698.0170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 697.8170 0.0000 698.0170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 697.8170 0.0000 698.0170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 697.8170 0.0000 698.0170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[125]

  PIN O[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 697.1340 0.0000 697.3340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 697.1340 0.0000 697.3340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 697.1340 0.0000 697.3340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 697.1340 0.0000 697.3340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 697.1340 0.0000 697.3340 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[124]

  PIN O[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 701.2380 0.0000 701.4380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 701.2380 0.0000 701.4380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 701.2380 0.0000 701.4380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 701.2380 0.0000 701.4380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 701.2380 0.0000 701.4380 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[127]

  PIN I[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 700.5530 0.0000 700.7530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 700.5530 0.0000 700.7530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 700.5530 0.0000 700.7530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 700.5530 0.0000 700.7530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 700.5530 0.0000 700.7530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[127]

  PIN O[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 699.8700 0.0000 700.0700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 699.8700 0.0000 700.0700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 699.8700 0.0000 700.0700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 699.8700 0.0000 700.0700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 699.8700 0.0000 700.0700 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[126]

  PIN I[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 699.1850 0.0000 699.3850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 699.1850 0.0000 699.3850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 699.1850 0.0000 699.3850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 699.1850 0.0000 699.3850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 699.1850 0.0000 699.3850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[126]

  PIN O[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 676.6140 0.0000 676.8140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 676.6140 0.0000 676.8140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 676.6140 0.0000 676.8140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 676.6140 0.0000 676.8140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 676.6140 0.0000 676.8140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[109]

  PIN O[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 675.2460 0.0000 675.4460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 675.2460 0.0000 675.4460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 675.2460 0.0000 675.4460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 675.2460 0.0000 675.4460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 675.2460 0.0000 675.4460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[108]

  PIN I[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 675.9290 0.0000 676.1290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 675.9290 0.0000 676.1290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 675.9290 0.0000 676.1290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 675.9290 0.0000 676.1290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 675.9290 0.0000 676.1290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[109]

  PIN O[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 680.7180 0.0000 680.9180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 680.7180 0.0000 680.9180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 680.7180 0.0000 680.9180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 680.7180 0.0000 680.9180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 680.7180 0.0000 680.9180 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[112]

  PIN O[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 679.3500 0.0000 679.5500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 679.3500 0.0000 679.5500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 679.3500 0.0000 679.5500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 679.3500 0.0000 679.5500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 679.3500 0.0000 679.5500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[111]

  PIN I[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 680.0330 0.0000 680.2330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 680.0330 0.0000 680.2330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 680.0330 0.0000 680.2330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 680.0330 0.0000 680.2330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 680.0330 0.0000 680.2330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[112]

  PIN I[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 678.6650 0.0000 678.8650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 678.6650 0.0000 678.8650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 678.6650 0.0000 678.8650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 678.6650 0.0000 678.8650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 678.6650 0.0000 678.8650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[111]

  PIN I[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 684.1370 0.0000 684.3370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 684.1370 0.0000 684.3370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 684.1370 0.0000 684.3370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 684.1370 0.0000 684.3370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 684.1370 0.0000 684.3370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[115]

  PIN O[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 683.4540 0.0000 683.6540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 683.4540 0.0000 683.6540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 683.4540 0.0000 683.6540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 683.4540 0.0000 683.6540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 683.4540 0.0000 683.6540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[114]

  PIN I[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 682.7690 0.0000 682.9690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 682.7690 0.0000 682.9690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 682.7690 0.0000 682.9690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 682.7690 0.0000 682.9690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 682.7690 0.0000 682.9690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[114]

  PIN I[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 681.4010 0.0000 681.6010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 681.4010 0.0000 681.6010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 681.4010 0.0000 681.6010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 681.4010 0.0000 681.6010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 681.4010 0.0000 681.6010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[113]

  PIN O[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 682.0860 0.0000 682.2860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 682.0860 0.0000 682.2860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 682.0860 0.0000 682.2860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 682.0860 0.0000 682.2860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 682.0860 0.0000 682.2860 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[113]

  PIN I[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 686.8730 0.0000 687.0730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 686.8730 0.0000 687.0730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 686.8730 0.0000 687.0730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 686.8730 0.0000 687.0730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 686.8730 0.0000 687.0730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[117]

  PIN O[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 686.1900 0.0000 686.3900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 686.1900 0.0000 686.3900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 686.1900 0.0000 686.3900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 686.1900 0.0000 686.3900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 686.1900 0.0000 686.3900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[116]

  PIN O[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 684.8220 0.0000 685.0220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 684.8220 0.0000 685.0220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 684.8220 0.0000 685.0220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 684.8220 0.0000 685.0220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 684.8220 0.0000 685.0220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[115]

  PIN I[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 685.5050 0.0000 685.7050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 685.5050 0.0000 685.7050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 685.5050 0.0000 685.7050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 685.5050 0.0000 685.7050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 685.5050 0.0000 685.7050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[116]

  PIN I[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 689.6090 0.0000 689.8090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 689.6090 0.0000 689.8090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 689.6090 0.0000 689.8090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 689.6090 0.0000 689.8090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 689.6090 0.0000 689.8090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[119]

  PIN O[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 690.2940 0.0000 690.4940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 690.2940 0.0000 690.4940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 690.2940 0.0000 690.4940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 690.2940 0.0000 690.4940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 690.2940 0.0000 690.4940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[119]

  PIN I[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 688.2410 0.0000 688.4410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 688.2410 0.0000 688.4410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 688.2410 0.0000 688.4410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 688.2410 0.0000 688.4410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 688.2410 0.0000 688.4410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[118]

  PIN I[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 663.6170 0.0000 663.8170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 663.6170 0.0000 663.8170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 663.6170 0.0000 663.8170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 663.6170 0.0000 663.8170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 663.6170 0.0000 663.8170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[100]

  PIN O[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 664.3020 0.0000 664.5020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 664.3020 0.0000 664.5020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 664.3020 0.0000 664.5020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 664.3020 0.0000 664.5020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 664.3020 0.0000 664.5020 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[100]

  PIN O[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 662.9340 0.0000 663.1340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 662.9340 0.0000 663.1340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 662.9340 0.0000 663.1340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 662.9340 0.0000 663.1340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 662.9340 0.0000 663.1340 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[99]

  PIN O[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 668.4060 0.0000 668.6060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 668.4060 0.0000 668.6060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 668.4060 0.0000 668.6060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 668.4060 0.0000 668.6060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 668.4060 0.0000 668.6060 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[103]

  PIN I[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 667.7210 0.0000 667.9210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 667.7210 0.0000 667.9210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 667.7210 0.0000 667.9210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 667.7210 0.0000 667.9210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 667.7210 0.0000 667.9210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[103]

  PIN I[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 666.3530 0.0000 666.5530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 666.3530 0.0000 666.5530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 666.3530 0.0000 666.5530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 666.3530 0.0000 666.5530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 666.3530 0.0000 666.5530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[102]

  PIN O[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 667.0380 0.0000 667.2380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 667.0380 0.0000 667.2380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 667.0380 0.0000 667.2380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 667.0380 0.0000 667.2380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 667.0380 0.0000 667.2380 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[102]

  PIN I[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 671.8250 0.0000 672.0250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 671.8250 0.0000 672.0250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 671.8250 0.0000 672.0250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 671.8250 0.0000 672.0250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 671.8250 0.0000 672.0250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[106]

  PIN O[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 671.1420 0.0000 671.3420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 671.1420 0.0000 671.3420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 671.1420 0.0000 671.3420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 671.1420 0.0000 671.3420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 671.1420 0.0000 671.3420 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[105]

  PIN O[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 669.7740 0.0000 669.9740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 669.7740 0.0000 669.9740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 669.7740 0.0000 669.9740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 669.7740 0.0000 669.9740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 669.7740 0.0000 669.9740 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[104]

  PIN I[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 670.4570 0.0000 670.6570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 670.4570 0.0000 670.6570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 670.4570 0.0000 670.6570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 670.4570 0.0000 670.6570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 670.4570 0.0000 670.6570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[105]

  PIN I[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 669.0890 0.0000 669.2890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 669.0890 0.0000 669.2890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 669.0890 0.0000 669.2890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 669.0890 0.0000 669.2890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 669.0890 0.0000 669.2890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[104]

  PIN I[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 674.5610 0.0000 674.7610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 674.5610 0.0000 674.7610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 674.5610 0.0000 674.7610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 674.5610 0.0000 674.7610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 674.5610 0.0000 674.7610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[108]

  PIN I[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 673.1930 0.0000 673.3930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 673.1930 0.0000 673.3930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 673.1930 0.0000 673.3930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 673.1930 0.0000 673.3930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 673.1930 0.0000 673.3930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[107]

  PIN O[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 673.8780 0.0000 674.0780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 673.8780 0.0000 674.0780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 673.8780 0.0000 674.0780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 673.8780 0.0000 674.0780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 673.8780 0.0000 674.0780 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[107]

  PIN O[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 672.5100 0.0000 672.7100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 672.5100 0.0000 672.7100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 672.5100 0.0000 672.7100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 672.5100 0.0000 672.7100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 672.5100 0.0000 672.7100 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[106]

  PIN O[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 677.9820 0.0000 678.1820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 677.9820 0.0000 678.1820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 677.9820 0.0000 678.1820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 677.9820 0.0000 678.1820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 677.9820 0.0000 678.1820 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[110]

  PIN I[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 677.2970 0.0000 677.4970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 677.2970 0.0000 677.4970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 677.2970 0.0000 677.4970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 677.2970 0.0000 677.4970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 677.2970 0.0000 677.4970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[110]

  PIN O[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 651.9900 0.0000 652.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 651.9900 0.0000 652.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 651.9900 0.0000 652.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 651.9900 0.0000 652.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 651.9900 0.0000 652.1900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[91]

  PIN I[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 651.3050 0.0000 651.5050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 651.3050 0.0000 651.5050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 651.3050 0.0000 651.5050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 651.3050 0.0000 651.5050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 651.3050 0.0000 651.5050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[91]

  PIN O[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 653.3580 0.0000 653.5580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 653.3580 0.0000 653.5580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 653.3580 0.0000 653.5580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 653.3580 0.0000 653.5580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 653.3580 0.0000 653.5580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[92]

  PIN I[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 652.6730 0.0000 652.8730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 652.6730 0.0000 652.8730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 652.6730 0.0000 652.8730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 652.6730 0.0000 652.8730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 652.6730 0.0000 652.8730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[92]

  PIN I[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 655.4090 0.0000 655.6090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 655.4090 0.0000 655.6090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 655.4090 0.0000 655.6090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 655.4090 0.0000 655.6090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 655.4090 0.0000 655.6090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[94]

  PIN O[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 656.0940 0.0000 656.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 656.0940 0.0000 656.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 656.0940 0.0000 656.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 656.0940 0.0000 656.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 656.0940 0.0000 656.2940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[94]

  PIN O[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 654.7260 0.0000 654.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 654.7260 0.0000 654.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 654.7260 0.0000 654.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 654.7260 0.0000 654.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 654.7260 0.0000 654.9260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[93]

  PIN I[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 654.0410 0.0010 654.2410 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 654.0410 0.0010 654.2410 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 654.0410 0.0000 654.2410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 654.0410 0.0000 654.2410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 654.0410 0.0000 654.2410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[93]

  PIN I[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 659.5130 0.0000 659.7130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 659.5130 0.0000 659.7130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 659.5130 0.0000 659.7130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 659.5130 0.0000 659.7130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 659.5130 0.0000 659.7130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[97]

  PIN O[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 658.8300 0.0000 659.0300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 658.8300 0.0000 659.0300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 658.8300 0.0000 659.0300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 658.8300 0.0000 659.0300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 658.8300 0.0000 659.0300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[96]

  PIN I[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 658.1450 0.0000 658.3450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 658.1450 0.0000 658.3450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 658.1450 0.0000 658.3450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 658.1450 0.0000 658.3450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 658.1450 0.0000 658.3450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[96]

  PIN O[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 657.4620 0.0000 657.6620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 657.4620 0.0000 657.6620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 657.4620 0.0000 657.6620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 657.4620 0.0000 657.6620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 657.4620 0.0000 657.6620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[95]

  PIN I[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 656.7770 0.0000 656.9770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 656.7770 0.0000 656.9770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 656.7770 0.0000 656.9770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 656.7770 0.0000 656.9770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 656.7770 0.0000 656.9770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[95]

  PIN I[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 662.2490 0.0000 662.4490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 662.2490 0.0000 662.4490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 662.2490 0.0000 662.4490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 662.2490 0.0000 662.4490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 662.2490 0.0000 662.4490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[99]

  PIN O[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 661.5660 0.0000 661.7660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 661.5660 0.0000 661.7660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 661.5660 0.0000 661.7660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 661.5660 0.0000 661.7660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 661.5660 0.0000 661.7660 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O[98]

  PIN I[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 660.8810 0.0000 661.0810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 660.8810 0.0000 661.0810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 660.8810 0.0000 661.0810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 660.8810 0.0000 661.0810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 660.8810 0.0000 661.0810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[98]
  OBS
    LAYER M2 ;
      RECT 0.0000 0.0000 526.1170 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 287.3560 722.2880 292.5510 ;
      RECT 0.0000 272.9260 723.1820 287.3560 ;
      RECT 0.0000 271.3260 722.2820 272.9260 ;
      RECT 721.6810 289.2990 723.1820 290.9510 ;
      RECT 0.0000 265.6960 723.1820 271.3260 ;
      RECT 0.0000 262.5060 722.2820 265.6960 ;
      RECT 0.0000 256.8760 723.1820 262.5060 ;
      RECT 0.0000 253.6860 722.2820 256.8760 ;
      RECT 0.0000 248.0600 723.1820 253.6860 ;
      RECT 0.0000 244.8700 722.2820 248.0600 ;
      RECT 0.0000 90.3700 723.1820 244.8700 ;
      RECT 0.0000 88.4090 722.2820 90.3700 ;
      RECT 0.0000 18.1900 723.1820 88.4090 ;
      RECT 0.0000 16.1280 722.2820 18.1900 ;
      RECT 0.0000 10.7200 723.1820 16.1280 ;
      RECT 0.0000 9.1200 722.2820 10.7200 ;
      RECT 0.0000 0.9000 723.1820 9.1200 ;
      RECT 0.0000 0.0000 526.1170 0.9000 ;
      RECT 702.8110 0.0000 723.1820 9.1200 ;
      RECT 702.8110 0.0000 723.1820 0.9000 ;
      RECT 0.0000 292.5510 723.1820 309.5940 ;
      RECT 0.0000 272.9260 722.2880 309.5940 ;
    LAYER M1 ;
      RECT 722.3820 246.3700 723.1820 246.5600 ;
      RECT 722.3820 255.1860 723.1820 255.3760 ;
      RECT 722.3820 264.0060 723.1820 264.1960 ;
      RECT 721.6810 289.1990 723.1820 291.0510 ;
      RECT 0.0000 265.5960 723.1820 271.4260 ;
      RECT 0.0000 262.6060 722.3820 265.5960 ;
      RECT 0.0000 256.7760 723.1820 262.6060 ;
      RECT 0.0000 253.7860 722.3820 256.7760 ;
      RECT 0.0000 247.9600 723.1820 253.7860 ;
      RECT 0.0000 244.9700 722.3820 247.9600 ;
      RECT 0.0000 90.2700 723.1820 244.9700 ;
      RECT 0.0000 88.5090 722.3820 90.2700 ;
      RECT 0.0000 18.0900 723.1820 88.5090 ;
      RECT 0.0000 16.2280 722.3820 18.0900 ;
      RECT 0.0000 10.6200 723.1820 16.2280 ;
      RECT 0.0000 9.2200 722.3820 10.6200 ;
      RECT 0.0000 0.8000 723.1820 9.2200 ;
      RECT 0.0000 0.0000 526.2170 0.8000 ;
      RECT 702.7110 0.0000 723.1820 9.2200 ;
      RECT 702.7110 0.0000 723.1820 0.8000 ;
      RECT 0.0000 292.4510 723.1820 309.5940 ;
      RECT 0.0000 272.8260 722.3880 309.5940 ;
      RECT 0.0000 0.0000 526.2170 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 0.8000 722.3820 309.5940 ;
      RECT 0.0000 287.4560 722.3880 292.4510 ;
      RECT 0.0000 272.8260 723.1820 287.4560 ;
      RECT 0.0000 271.4260 722.3820 272.8260 ;
    LAYER PO ;
      RECT 0.0000 0.0000 723.1820 309.5940 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 723.1820 309.5940 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 723.1820 309.5940 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 723.1820 309.5940 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 723.1820 309.5940 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 723.1820 309.5940 ;
    LAYER M5 ;
      RECT 722.3510 308.5940 723.1820 309.5940 ;
      RECT 721.6810 289.2990 723.1820 290.9510 ;
      RECT 702.8110 0.0000 723.1820 0.9000 ;
      RECT 0.0000 0.0000 526.1170 0.9000 ;
      RECT 0.0000 265.6960 723.1820 271.3260 ;
      RECT 0.0000 262.5060 722.2820 265.6960 ;
      RECT 0.0000 256.8760 723.1820 262.5060 ;
      RECT 0.0000 253.6860 722.2820 256.8760 ;
      RECT 0.0000 248.0600 723.1820 253.6860 ;
      RECT 0.0000 244.8700 722.2820 248.0600 ;
      RECT 0.0000 90.3700 723.1820 244.8700 ;
      RECT 0.0000 88.4090 722.2820 90.3700 ;
      RECT 0.0000 18.1900 723.1820 88.4090 ;
      RECT 0.0000 16.1280 722.2820 18.1900 ;
      RECT 0.0000 10.7200 723.1820 16.1280 ;
      RECT 0.0000 9.1200 722.2820 10.7200 ;
      RECT 0.0000 0.9010 723.1820 9.1200 ;
      RECT 0.0000 0.9000 527.4850 0.9010 ;
      RECT 529.0850 0.9000 590.4130 0.9010 ;
      RECT 592.0130 0.9000 653.3410 0.9010 ;
      RECT 654.9410 0.9000 723.1820 9.1200 ;
      RECT 654.9410 0.9000 723.1820 0.9010 ;
      RECT 0.0000 0.9000 527.4850 308.5940 ;
      RECT 0.0000 292.5510 723.1820 308.5940 ;
      RECT 0.0000 272.9260 722.2880 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 0.9010 722.2820 308.5940 ;
      RECT 0.0000 287.3560 722.2880 292.5510 ;
      RECT 0.0000 272.9260 723.1820 287.3560 ;
      RECT 0.0000 271.3260 722.2820 272.9260 ;
      RECT 529.0850 0.9000 590.4130 308.5940 ;
      RECT 592.0130 0.9000 653.3410 308.5940 ;
    LAYER M4 ;
      RECT 721.6810 289.2990 723.1820 290.9510 ;
      RECT 702.8110 0.0000 723.1820 0.9000 ;
      RECT 0.0000 0.0000 526.1170 0.9000 ;
      RECT 0.0000 265.6960 723.1820 271.3260 ;
      RECT 0.0000 262.5060 722.2820 265.6960 ;
      RECT 0.0000 256.8760 723.1820 262.5060 ;
      RECT 0.0000 253.6860 722.2820 256.8760 ;
      RECT 0.0000 248.0600 723.1820 253.6860 ;
      RECT 0.0000 244.8700 722.2820 248.0600 ;
      RECT 0.0000 90.3700 723.1820 244.8700 ;
      RECT 0.0000 88.4090 722.2820 90.3700 ;
      RECT 0.0000 18.1900 723.1820 88.4090 ;
      RECT 0.0000 16.1280 722.2820 18.1900 ;
      RECT 0.0000 10.7200 723.1820 16.1280 ;
      RECT 0.0000 9.1200 722.2820 10.7200 ;
      RECT 0.0000 0.9010 723.1820 9.1200 ;
      RECT 0.0000 0.9000 527.4850 0.9010 ;
      RECT 529.0850 0.9000 590.4130 0.9010 ;
      RECT 592.0130 0.9000 653.3410 0.9010 ;
      RECT 654.9410 0.9000 723.1820 9.1200 ;
      RECT 654.9410 0.9000 723.1820 0.9010 ;
      RECT 0.0000 0.9000 527.4850 309.5940 ;
      RECT 0.0000 292.5510 723.1820 309.5940 ;
      RECT 0.0000 272.9260 722.2880 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 0.9010 722.2820 309.5940 ;
      RECT 0.0000 287.3560 722.2880 292.5510 ;
      RECT 0.0000 272.9260 723.1820 287.3560 ;
      RECT 0.0000 271.3260 722.2820 272.9260 ;
      RECT 529.0850 0.9000 590.4130 309.5940 ;
      RECT 592.0130 0.9000 653.3410 309.5940 ;
    LAYER M3 ;
      RECT 721.6810 289.2990 723.1820 290.9510 ;
      RECT 0.0000 265.6960 723.1820 271.3260 ;
      RECT 0.0000 262.5060 722.2820 265.6960 ;
      RECT 0.0000 256.8760 723.1820 262.5060 ;
      RECT 0.0000 253.6860 722.2820 256.8760 ;
      RECT 0.0000 248.0600 723.1820 253.6860 ;
      RECT 0.0000 244.8700 722.2820 248.0600 ;
      RECT 0.0000 90.3700 723.1820 244.8700 ;
      RECT 0.0000 88.4090 722.2820 90.3700 ;
      RECT 0.0000 18.1900 723.1820 88.4090 ;
      RECT 0.0000 16.1280 722.2820 18.1900 ;
      RECT 0.0000 10.7200 723.1820 16.1280 ;
      RECT 0.0000 9.1200 722.2820 10.7200 ;
      RECT 0.0000 0.9000 723.1820 9.1200 ;
      RECT 0.0000 0.0000 526.1170 0.9000 ;
      RECT 702.8110 0.0000 723.1820 9.1200 ;
      RECT 702.8110 0.0000 723.1820 0.9000 ;
      RECT 0.0000 292.5510 723.1820 309.5940 ;
      RECT 0.0000 272.9260 722.2880 309.5940 ;
      RECT 0.0000 0.0000 526.1170 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 0.9000 722.2820 309.5940 ;
      RECT 0.0000 287.3560 722.2880 292.5510 ;
      RECT 0.0000 272.9260 723.1820 287.3560 ;
      RECT 0.0000 271.3260 722.2820 272.9260 ;
  END
END SRAMLP1RW512x128

MACRO SRAMLP1RW1024x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 110.903 BY 244.693 ;
  SYMMETRY X Y R90 ;

  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 36.4940 110.9030 36.6940 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 36.4940 110.9030 36.6940 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 36.4940 110.9030 36.6940 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 36.4940 110.9030 36.6940 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 36.4940 110.9030 36.6940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[9]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.5740 0.0000 86.7740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.5740 0.0000 86.7740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.5740 0.0000 86.7740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.5740 0.0000 86.7740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.5740 0.0000 86.7740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.9200 0.0000 86.1200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.9200 0.0000 86.1200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.9200 0.0000 86.1200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.9200 0.0000 86.1200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.9200 0.0000 86.1200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[7]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.2060 0.0000 85.4060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.2060 0.0000 85.4060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.2060 0.0000 85.4060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.2060 0.0000 85.4060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.2060 0.0000 85.4060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 41.2170 110.9030 41.4170 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 41.2170 110.9030 41.4170 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 41.2170 110.9030 41.4170 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 41.2170 110.9030 41.4170 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 41.2170 110.9030 41.4170 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[7]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.6970 16.8900 110.8940 17.0900 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.6970 16.8900 110.8940 17.0900 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.6970 16.8900 110.8940 17.0900 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.6970 16.8900 110.8940 17.0900 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.6970 16.8900 110.8940 17.0900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 9.8900 110.9030 10.0900 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 9.8900 110.9030 10.0900 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 9.8900 110.9030 10.0900 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 9.8900 110.9030 10.0900 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 9.8900 110.9030 10.0900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 198.4770 110.9030 198.6770 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 198.4770 110.9030 198.6770 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 198.4770 110.9030 198.6770 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 198.4770 110.9030 198.6770 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 198.4770 110.9030 198.6770 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 234.4560 110.9030 234.6560 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 234.4560 110.9030 234.6560 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 234.4560 110.9030 234.6560 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 234.4560 110.9030 234.6560 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 234.4560 110.9030 234.6560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 2.3360 244.3930 2.6350 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2340 244.3930 3.5340 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1340 244.3930 85.4340 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0340 244.3930 86.3350 244.6930 ;
    END
  END VDDL

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.6730 207.4910 110.8730 207.6910 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.6730 207.4910 110.8730 207.6910 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.6730 207.4910 110.8730 207.6910 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.6730 207.4910 110.8730 207.6910 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.6730 207.4910 110.8730 207.6910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 234.8690 110.9030 235.0690 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 234.8690 110.9030 235.0690 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 234.8690 110.9030 235.0690 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 234.8690 110.9030 235.0690 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 234.8690 110.9030 235.0690 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 237.9520 110.9030 238.1520 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 237.9520 110.9030 238.1520 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 237.9520 110.9030 238.1520 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 237.9520 110.9030 238.1520 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 237.9520 110.9030 238.1520 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 200.0670 110.9030 200.2670 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 200.0670 110.9030 200.2670 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 200.0670 110.9030 200.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 200.0670 110.9030 200.2670 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 200.0670 110.9030 200.2670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.4500 0.0000 80.6500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.4500 0.0000 80.6500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.4500 0.0000 80.6500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.4500 0.0000 80.6500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.4500 0.0000 80.6500 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278508 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278508 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[3]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.7340 0.0000 79.9340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.7340 0.0000 79.9340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.7340 0.0000 79.9340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.7340 0.0000 79.9340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.7340 0.0000 79.9340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.6260 189.6490 110.8260 189.8490 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.6260 189.6490 110.8260 189.8490 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.6260 189.6490 110.8260 189.8490 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.6260 189.6490 110.8260 189.8490 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.6260 189.6490 110.8260 189.8490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 182.4180 110.9030 182.6180 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 182.4180 110.9030 182.6180 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 182.4180 110.9030 182.6180 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 182.4180 110.9030 182.6180 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 182.4180 110.9030 182.6180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 180.8420 110.9030 181.0420 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 180.8420 110.9030 181.0420 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 180.8420 110.9030 181.0420 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 180.8420 110.9030 181.0420 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 180.8420 110.9030 181.0420 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[6]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7020 17.3590 110.8990 17.5590 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7020 17.3590 110.8990 17.5590 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7020 17.3590 110.8990 17.5590 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7020 17.3590 110.8990 17.5590 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7020 17.3590 110.8990 17.5590 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7030 38.7700 110.9030 38.9700 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7030 38.7700 110.9030 38.9700 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7030 38.7700 110.9030 38.9700 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7030 38.7700 110.9030 38.9700 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7030 38.7700 110.9030 38.9700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[8]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.1730 0.0000 83.3730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.1730 0.0000 83.3730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.1730 0.0000 83.3730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.1730 0.0000 83.3730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.1730 0.0000 83.3730 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[5]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.6980 0.0000 77.8980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.6980 0.0000 77.8980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.6980 0.0000 77.8980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.6980 0.0000 77.8980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.6980 0.0000 77.8980 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[1]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.8040 0.0000 82.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.8040 0.0000 82.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.8040 0.0000 82.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.8040 0.0000 82.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.8040 0.0000 82.0040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[4]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.5430 0.0000 84.7430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.5430 0.0000 84.7430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.5430 0.0000 84.7430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.5430 0.0000 84.7430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.5430 0.0000 84.7430 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[6]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.3660 0.0000 78.5660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.3660 0.0000 78.5660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.3660 0.0000 78.5660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.3660 0.0000 78.5660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.3660 0.0000 78.5660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.4700 0.0000 82.6700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.4700 0.0000 82.6700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.4700 0.0000 82.6700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.4700 0.0000 82.6700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.4700 0.0000 82.6700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.1020 0.0000 81.3020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.1020 0.0000 81.3020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.1020 0.0000 81.3020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.1020 0.0000 81.3020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.1020 0.0000 81.3020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.0680 0.0000 79.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.0680 0.0000 79.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.0680 0.0000 79.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.0680 0.0000 79.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.0680 0.0000 79.2680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[2]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.0490 0.0000 89.2490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.0490 0.0000 89.2490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.0490 0.0000 89.2490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.0490 0.0000 89.2490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.0490 0.0000 89.2490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.6260 191.2390 110.8260 191.4390 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.6260 191.2390 110.8260 191.4390 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.6260 191.2390 110.8260 191.4390 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.6260 191.2390 110.8260 191.4390 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.6260 191.2390 110.8260 191.4390 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.3280 0.0000 76.5280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.3280 0.0000 76.5280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.3280 0.0000 76.5280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.3280 0.0000 76.5280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.3280 0.0000 76.5280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.27238 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27238 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[0]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.8380 0.0000 84.0380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.8380 0.0000 84.0380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.8380 0.0000 84.0380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.8380 0.0000 84.0380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.8380 0.0000 84.0380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.9980 0.0000 77.1980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.9980 0.0000 77.1980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.9980 0.0000 77.1980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.9980 0.0000 77.1980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.9980 0.0000 77.1980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 1.4330 244.3930 1.7340 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.8350 244.3930 88.1350 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.5350 244.3930 0.8340 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.9350 244.3930 87.2340 244.6930 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 1.8850 244.3930 2.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.3850 244.3930 6.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6830 244.3930 3.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7850 244.3930 3.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.5860 244.3930 4.8850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.4840 244.3930 5.7840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0840 244.3930 0.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.8850 244.3930 11.1840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.2850 244.3930 7.5850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.0840 244.3930 9.3850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.1840 244.3930 8.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.9850 244.3930 10.2840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.4850 244.3930 14.7840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6840 244.3930 12.9850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7840 244.3930 12.0840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.5840 244.3930 13.8850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.2840 244.3930 16.5840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.3850 244.3930 15.6840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.9850 244.3930 19.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0840 244.3930 18.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1850 244.3930 17.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.8840 244.3930 20.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.7850 244.3930 21.0840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.4850 244.3930 23.7850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.1860 244.3930 26.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.3850 244.3930 24.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.2830 244.3930 25.5840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.5840 244.3930 22.8850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.6840 244.3930 21.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.0840 244.3930 27.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.8850 244.3930 29.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.6840 244.3930 30.9850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.7840 244.3930 30.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.9850 244.3930 28.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.2840 244.3930 34.5850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.4850 244.3930 32.7840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.3840 244.3930 33.6840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.1840 244.3930 35.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.5850 244.3930 31.8840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.0850 244.3930 36.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.5850 244.3930 40.8850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.6840 244.3930 39.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.7850 244.3930 39.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.8840 244.3930 38.1840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.9850 244.3930 37.2840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.0850 244.3930 45.3850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.4840 244.3930 41.7850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.1840 244.3930 44.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.3850 244.3930 42.6840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.2840 244.3930 43.5840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.6840 244.3930 48.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.7860 244.3930 48.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.9850 244.3930 46.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.8830 244.3930 47.1840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.5850 244.3930 49.8850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.0850 244.3930 54.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.9840 244.3930 55.2840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.4850 244.3930 50.7850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.2840 244.3930 52.5850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.3840 244.3930 51.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.1850 244.3930 53.4840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.6850 244.3930 57.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.8840 244.3930 56.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.7840 244.3930 57.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.4840 244.3930 59.7840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.5850 244.3930 58.8840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.1850 244.3930 62.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.2840 244.3930 61.5840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.3850 244.3930 60.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.0840 244.3930 63.3850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.9850 244.3930 64.2840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.8840 244.3930 65.1840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.3860 244.3930 69.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.5850 244.3930 67.8850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.4830 244.3930 68.7840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.7840 244.3930 66.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.6850 244.3930 66.9850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.2840 244.3930 70.5840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.0850 244.3930 72.3850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.8840 244.3930 74.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.9840 244.3930 73.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.1850 244.3930 71.4850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.2850 244.3930 79.5840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.4840 244.3930 77.7850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.6850 244.3930 75.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.5840 244.3930 76.8840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.3840 244.3930 78.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.7850 244.3930 75.0840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.7850 244.3930 84.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.8840 244.3930 83.1840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.9850 244.3930 82.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.0840 244.3930 81.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.1850 244.3930 80.4840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.2850 244.3930 88.5850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.6840 244.3930 84.9850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.3840 244.3930 87.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.5850 244.3930 85.8840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.4840 244.3930 86.7840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.1840 244.3930 89.4840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.9840 244.3930 91.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.8840 244.3930 92.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.7840 244.3930 93.0850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.6850 244.3930 93.9850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.0840 244.3930 90.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.1850 244.3930 98.4840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.5850 244.3930 94.8840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.4850 244.3930 95.7850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.3840 244.3930 96.6840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.2850 244.3930 97.5850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.9840 244.3930 100.2850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.8840 244.3930 101.1850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.0840 244.3930 99.3840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.7850 244.3930 102.0840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.6850 244.3930 102.9840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.4840 244.3930 104.7850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.3840 244.3930 105.6850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.2850 244.3930 106.5850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.1840 244.3930 107.4840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.0850 244.3930 108.3850 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.5840 244.3930 103.8840 244.6930 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.9840 244.3930 1.2850 244.6930 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0000 37.2940 110.1030 180.2420 ;
      RECT 0.0000 40.6170 110.1030 42.0170 ;
      RECT 0.0000 39.5700 110.1030 40.6170 ;
      RECT 0.0000 38.1700 110.1030 39.5700 ;
      RECT 0.0000 37.2940 110.1030 38.1700 ;
      RECT 89.8490 0.0000 110.9030 0.8000 ;
      RECT 0.0000 0.0000 75.7280 0.8000 ;
      RECT 0.0000 0.0000 75.7280 9.2900 ;
      RECT 0.0000 0.8000 110.9030 9.2900 ;
      RECT 89.8490 0.0000 110.9030 9.2900 ;
      RECT 0.0000 35.8940 110.1030 180.2420 ;
      RECT 0.0000 35.8940 110.1030 180.2420 ;
      RECT 0.0000 35.8940 110.1030 180.2420 ;
      RECT 0.0000 35.8940 110.1030 180.2420 ;
      RECT 0.0000 35.8940 110.1030 180.2420 ;
      RECT 0.0000 35.8940 110.1030 180.2420 ;
      RECT 0.0000 35.8940 110.1030 42.0170 ;
      RECT 0.0000 35.8940 110.1030 42.0170 ;
      RECT 0.0000 35.8940 110.1030 40.6170 ;
      RECT 0.0000 35.8940 110.1030 40.6170 ;
      RECT 0.0000 35.8940 110.1030 40.6170 ;
      RECT 0.0000 35.8940 110.1030 40.6170 ;
      RECT 0.0000 35.8940 110.1030 40.6170 ;
      RECT 0.0000 35.8940 110.1030 40.6170 ;
      RECT 0.0000 35.8940 110.1030 37.2940 ;
      RECT 0.0000 18.1590 110.9030 35.8940 ;
      RECT 0.0000 17.6900 110.1020 35.8940 ;
      RECT 0.0000 17.6900 110.1020 35.8940 ;
      RECT 0.0000 17.6900 110.1020 18.1590 ;
      RECT 0.0000 16.2900 110.0970 17.6900 ;
      RECT 0.0000 10.6900 110.0970 17.6900 ;
      RECT 0.0000 10.6900 110.0970 17.6900 ;
      RECT 0.0000 10.6900 110.9030 16.2900 ;
      RECT 0.0000 9.2900 110.1030 16.2900 ;
      RECT 0.0000 9.2900 110.1030 10.6900 ;
      RECT 110.0260 190.4490 110.9030 190.6390 ;
      RECT 110.1030 199.2770 110.9030 199.4670 ;
      RECT 110.1030 181.6420 110.9030 181.8180 ;
      RECT 110.1030 37.2940 110.9030 38.1700 ;
      RECT 110.1030 39.5700 110.9030 40.6170 ;
      RECT 87.3740 0.0000 88.4490 0.8000 ;
      RECT 109.4020 235.6690 110.9030 237.3520 ;
      RECT 0.0000 238.7520 110.9030 244.6930 ;
      RECT 0.0000 237.3520 110.1030 238.7520 ;
      RECT 0.0000 235.6690 110.1030 238.7520 ;
      RECT 0.0000 235.6690 110.1030 237.3520 ;
      RECT 0.0000 233.8560 110.1030 244.6930 ;
      RECT 0.0000 233.8560 110.1030 244.6930 ;
      RECT 0.0000 233.8560 110.1030 244.6930 ;
      RECT 0.0000 233.8560 110.1030 244.6930 ;
      RECT 0.0000 233.8560 110.1030 238.7520 ;
      RECT 0.0000 233.8560 110.1030 237.3520 ;
      RECT 0.0000 233.8560 110.1030 237.3520 ;
      RECT 0.0000 233.8560 110.1030 237.3520 ;
      RECT 0.0000 233.8560 110.1030 235.6690 ;
      RECT 0.0000 208.2910 110.9030 233.8560 ;
      RECT 0.0000 206.8910 110.0730 233.8560 ;
      RECT 0.0000 206.8910 110.0730 208.2910 ;
      RECT 0.0000 200.8670 110.9030 206.8910 ;
      RECT 0.0000 199.4670 110.1030 200.8670 ;
      RECT 0.0000 199.2770 110.1030 199.4670 ;
      RECT 0.0000 192.0390 110.1030 206.8910 ;
      RECT 0.0000 192.0390 110.1030 206.8910 ;
      RECT 0.0000 192.0390 110.1030 206.8910 ;
      RECT 0.0000 192.0390 110.1030 206.8910 ;
      RECT 0.0000 192.0390 110.1030 206.8910 ;
      RECT 0.0000 192.0390 110.1030 206.8910 ;
      RECT 0.0000 192.0390 110.1030 199.4670 ;
      RECT 0.0000 192.0390 110.1030 199.4670 ;
      RECT 0.0000 192.0390 110.1030 199.4670 ;
      RECT 0.0000 197.8770 110.1030 199.2770 ;
      RECT 0.0000 192.0390 110.9030 197.8770 ;
      RECT 0.0000 190.4490 110.0260 197.8770 ;
      RECT 0.0000 190.4490 110.0260 197.8770 ;
      RECT 0.0000 190.4490 110.0260 197.8770 ;
      RECT 0.0000 190.6390 110.0260 192.0390 ;
      RECT 0.0000 190.4490 110.0260 190.6390 ;
      RECT 0.0000 189.0490 110.0260 197.8770 ;
      RECT 0.0000 189.0490 110.0260 197.8770 ;
      RECT 0.0000 189.0490 110.0260 197.8770 ;
      RECT 0.0000 189.0490 110.0260 190.4490 ;
      RECT 0.0000 183.2180 110.9030 189.0490 ;
      RECT 0.0000 181.6420 110.1030 189.0490 ;
      RECT 0.0000 181.6420 110.1030 189.0490 ;
      RECT 0.0000 181.6420 110.1030 189.0490 ;
      RECT 0.0000 181.8180 110.1030 183.2180 ;
      RECT 0.0000 181.6420 110.1030 181.8180 ;
      RECT 0.0000 180.2420 110.1030 189.0490 ;
      RECT 0.0000 180.2420 110.1030 189.0490 ;
      RECT 0.0000 180.2420 110.1030 189.0490 ;
      RECT 0.0000 180.2420 110.1030 181.6420 ;
      RECT 0.0000 42.0170 110.9030 180.2420 ;
      RECT 0.0000 38.1700 110.1030 180.2420 ;
      RECT 0.0000 38.1700 110.1030 180.2420 ;
    LAYER PO ;
      RECT 0.0000 0.0000 110.9030 244.6930 ;
    LAYER M3 ;
      RECT 0.0000 0.9000 110.9030 9.1900 ;
      RECT 0.0000 0.0000 75.6280 0.9000 ;
      RECT 89.9490 0.0000 110.9030 9.1900 ;
      RECT 89.9490 0.0000 110.9030 0.9000 ;
      RECT 0.0000 200.9670 110.9030 206.7910 ;
      RECT 0.0000 192.1390 110.0030 206.7910 ;
      RECT 0.0000 197.7770 110.0030 200.9670 ;
      RECT 0.0000 192.1390 110.9030 197.7770 ;
      RECT 0.0000 188.9490 109.9260 192.1390 ;
      RECT 0.0000 0.9000 109.9260 192.1390 ;
      RECT 0.0000 238.8520 110.9030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 192.1390 109.9730 244.6930 ;
      RECT 0.0000 0.0000 75.6280 244.6930 ;
      RECT 0.0000 237.2520 110.0030 238.8520 ;
      RECT 0.0000 235.7690 110.0030 237.2520 ;
      RECT 0.0000 233.7560 110.0030 235.7690 ;
      RECT 0.0000 208.3910 110.9030 233.7560 ;
      RECT 0.0000 206.7910 109.9730 208.3910 ;
      RECT 87.4740 0.0000 88.3490 0.9000 ;
      RECT 110.0030 235.7690 110.9030 237.2520 ;
      RECT 110.0030 37.3940 110.9030 38.0700 ;
      RECT 110.0030 39.6700 110.9030 40.5170 ;
      RECT 0.0000 183.3180 110.9030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 17.7900 110.0020 188.9490 ;
      RECT 0.0000 0.9000 109.9970 188.9490 ;
      RECT 0.0000 180.1420 110.0030 183.3180 ;
      RECT 0.0000 42.1170 110.9030 180.1420 ;
      RECT 0.0000 40.5170 110.0030 42.1170 ;
      RECT 0.0000 39.6700 110.0030 40.5170 ;
      RECT 0.0000 38.0700 110.0030 39.6700 ;
      RECT 0.0000 37.3940 110.0030 38.0700 ;
      RECT 0.0000 35.7940 110.0030 37.3940 ;
      RECT 0.0000 18.2590 110.9030 35.7940 ;
      RECT 0.0000 17.7900 110.0020 18.2590 ;
      RECT 0.0000 16.1900 109.9970 17.7900 ;
      RECT 0.0000 10.7900 110.9030 16.1900 ;
      RECT 0.0000 0.9000 110.0030 16.1900 ;
      RECT 0.0000 9.1900 110.0030 10.7900 ;
    LAYER M2 ;
      RECT 110.0030 39.6700 110.9030 40.5170 ;
      RECT 110.0030 37.3940 110.9030 38.0700 ;
      RECT 110.0030 235.7690 110.9030 237.2520 ;
      RECT 87.4740 0.0000 88.3490 0.9000 ;
      RECT 0.0000 183.3180 110.9030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 17.7900 110.0020 188.9490 ;
      RECT 0.0000 0.9000 109.9970 188.9490 ;
      RECT 0.0000 180.1420 110.0030 183.3180 ;
      RECT 0.0000 42.1170 110.9030 180.1420 ;
      RECT 0.0000 40.5170 110.0030 42.1170 ;
      RECT 0.0000 39.6700 110.0030 40.5170 ;
      RECT 0.0000 38.0700 110.0030 39.6700 ;
      RECT 0.0000 37.3940 110.0030 38.0700 ;
      RECT 0.0000 35.7940 110.0030 37.3940 ;
      RECT 0.0000 18.2590 110.9030 35.7940 ;
      RECT 0.0000 17.7900 110.0020 18.2590 ;
      RECT 0.0000 16.1900 109.9970 17.7900 ;
      RECT 0.0000 10.7900 110.9030 16.1900 ;
      RECT 0.0000 0.9000 110.0030 16.1900 ;
      RECT 0.0000 9.1900 110.0030 10.7900 ;
      RECT 0.0000 0.9000 110.9030 9.1900 ;
      RECT 0.0000 0.0000 75.6280 0.9000 ;
      RECT 89.9490 0.0000 110.9030 9.1900 ;
      RECT 89.9490 0.0000 110.9030 0.9000 ;
      RECT 0.0000 200.9670 110.9030 206.7910 ;
      RECT 0.0000 192.1390 110.0030 206.7910 ;
      RECT 0.0000 197.7770 110.0030 200.9670 ;
      RECT 0.0000 192.1390 110.9030 197.7770 ;
      RECT 0.0000 188.9490 109.9260 192.1390 ;
      RECT 0.0000 0.9000 109.9260 192.1390 ;
      RECT 0.0000 238.8520 110.9030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 192.1390 109.9730 244.6930 ;
      RECT 0.0000 0.0000 75.6280 244.6930 ;
      RECT 0.0000 237.2520 110.0030 238.8520 ;
      RECT 0.0000 235.7690 110.0030 237.2520 ;
      RECT 0.0000 233.7560 110.0030 235.7690 ;
      RECT 0.0000 208.3910 110.9030 233.7560 ;
      RECT 0.0000 206.7910 109.9730 208.3910 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 110.9030 244.6930 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 110.9030 244.6930 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 110.9030 244.6930 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 110.9030 244.6930 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 110.9030 244.6930 ;
    LAYER M5 ;
      RECT 87.4740 0.0000 88.3490 0.9000 ;
      RECT 109.0850 243.6930 110.9030 244.6930 ;
      RECT 109.0850 243.1920 110.9030 244.6930 ;
      RECT 110.0030 235.7690 110.9030 237.2520 ;
      RECT 110.0030 37.3940 110.9030 38.0700 ;
      RECT 110.0030 39.6700 110.9030 40.5170 ;
      RECT 0.0000 183.3180 110.9030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 17.7900 110.0020 188.9490 ;
      RECT 0.0000 0.9000 109.9970 188.9490 ;
      RECT 0.0000 180.1420 110.0030 183.3180 ;
      RECT 0.0000 42.1170 110.9030 180.1420 ;
      RECT 0.0000 40.5170 110.0030 42.1170 ;
      RECT 0.0000 39.6700 110.0030 40.5170 ;
      RECT 0.0000 38.0700 110.0030 39.6700 ;
      RECT 0.0000 37.3940 110.0030 38.0700 ;
      RECT 0.0000 35.7940 110.0030 37.3940 ;
      RECT 0.0000 18.2590 110.9030 35.7940 ;
      RECT 0.0000 17.7900 110.0020 18.2590 ;
      RECT 0.0000 16.1900 109.9970 17.7900 ;
      RECT 0.0000 10.7900 110.9030 16.1900 ;
      RECT 0.0000 0.9000 110.0030 16.1900 ;
      RECT 0.0000 9.1900 110.0030 10.7900 ;
      RECT 0.0000 0.9000 110.9030 9.1900 ;
      RECT 0.0000 0.0000 75.6280 0.9000 ;
      RECT 89.9490 0.0000 110.9030 9.1900 ;
      RECT 89.9490 0.0000 110.9030 0.9000 ;
      RECT 0.0000 200.9670 110.9030 206.7910 ;
      RECT 0.0000 192.1390 110.0030 206.7910 ;
      RECT 0.0000 197.7770 110.0030 200.9670 ;
      RECT 0.0000 192.1390 110.9030 197.7770 ;
      RECT 0.0000 188.9490 109.9260 192.1390 ;
      RECT 0.0000 0.9000 109.9260 192.1390 ;
      RECT 0.0000 238.8520 110.9030 243.6930 ;
      RECT 0.0000 208.3910 110.0030 243.6930 ;
      RECT 0.0000 208.3910 110.0030 243.6930 ;
      RECT 0.0000 208.3910 110.0030 243.6930 ;
      RECT 0.0000 192.1390 109.9730 243.6930 ;
      RECT 0.0000 0.0000 75.6280 243.6930 ;
      RECT 0.0000 237.2520 110.0030 238.8520 ;
      RECT 0.0000 235.7690 110.0030 237.2520 ;
      RECT 0.0000 233.7560 110.0030 235.7690 ;
      RECT 0.0000 208.3910 110.9030 233.7560 ;
      RECT 0.0000 206.7910 109.9730 208.3910 ;
    LAYER M4 ;
      RECT 87.4740 0.0000 88.3490 0.9000 ;
      RECT 110.0030 235.7690 110.9030 237.2520 ;
      RECT 110.0030 37.3940 110.9030 38.0700 ;
      RECT 110.0030 39.6700 110.9030 40.5170 ;
      RECT 0.0000 183.3180 110.9030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 18.2590 110.0030 188.9490 ;
      RECT 0.0000 17.7900 110.0020 188.9490 ;
      RECT 0.0000 0.9000 109.9970 188.9490 ;
      RECT 0.0000 180.1420 110.0030 183.3180 ;
      RECT 0.0000 42.1170 110.9030 180.1420 ;
      RECT 0.0000 40.5170 110.0030 42.1170 ;
      RECT 0.0000 39.6700 110.0030 40.5170 ;
      RECT 0.0000 38.0700 110.0030 39.6700 ;
      RECT 0.0000 37.3940 110.0030 38.0700 ;
      RECT 0.0000 35.7940 110.0030 37.3940 ;
      RECT 0.0000 18.2590 110.9030 35.7940 ;
      RECT 0.0000 17.7900 110.0020 18.2590 ;
      RECT 0.0000 16.1900 109.9970 17.7900 ;
      RECT 0.0000 10.7900 110.9030 16.1900 ;
      RECT 0.0000 0.9000 110.0030 16.1900 ;
      RECT 0.0000 9.1900 110.0030 10.7900 ;
      RECT 0.0000 0.9000 110.9030 9.1900 ;
      RECT 0.0000 0.0000 75.6280 0.9000 ;
      RECT 89.9490 0.0000 110.9030 9.1900 ;
      RECT 89.9490 0.0000 110.9030 0.9000 ;
      RECT 0.0000 200.9670 110.9030 206.7910 ;
      RECT 0.0000 192.1390 110.0030 206.7910 ;
      RECT 0.0000 197.7770 110.0030 200.9670 ;
      RECT 0.0000 192.1390 110.9030 197.7770 ;
      RECT 0.0000 188.9490 109.9260 192.1390 ;
      RECT 0.0000 0.9000 109.9260 192.1390 ;
      RECT 0.0000 238.8520 110.9030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 208.3910 110.0030 244.6930 ;
      RECT 0.0000 192.1390 109.9730 244.6930 ;
      RECT 0.0000 0.0000 75.6280 244.6930 ;
      RECT 0.0000 237.2520 110.0030 238.8520 ;
      RECT 0.0000 235.7690 110.0030 237.2520 ;
      RECT 0.0000 233.7560 110.0030 235.7690 ;
      RECT 0.0000 208.3910 110.9030 233.7560 ;
      RECT 0.0000 206.7910 109.9730 208.3910 ;
  END
END SRAMLP1RW1024x8

MACRO SRAMLP2RW16x4
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 55.645 BY 52.479 ;
  SYMMETRY X Y R90 ;

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.123568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.123568 LAYER M3 ;
    ANTENNAMAXAREACAR 33.06199 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.20189 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.34151 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAGATEAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.171326 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.171326 LAYER M2 ;
    ANTENNAMAXAREACAR 63.68736 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 70.90221 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 78.11658 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 85.33047 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[3]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.111148 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.111148 LAYER M3 ;
    ANTENNAMAXAREACAR 32.72265 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.86256 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.00221 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.111148 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.111148 LAYER M3 ;
    ANTENNAMAXAREACAR 32.72265 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.86256 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.00221 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[2]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.111148 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.111148 LAYER M3 ;
    ANTENNAMAXAREACAR 32.72265 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.86256 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.00221 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[0]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.42508 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.42508 LAYER M4 ;
    ANTENNAMAXAREACAR 14.04121 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.18236 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 17.2520 55.6450 17.4520 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 17.2520 55.6450 17.4520 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 17.2520 55.6450 17.4520 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 17.2520 55.6450 17.4520 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 17.2520 55.6450 17.4520 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0894 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.32626 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.32626 LAYER M4 ;
    ANTENNAMAXAREACAR 6.863049 LAYER M4 ;
    ANTENNAGATEAREA 0.0894 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.558346 LAYER M5 ;
    ANTENNAGATEAREA 0.0894 LAYER M6 ;
    ANTENNAGATEAREA 0.0894 LAYER M7 ;
    ANTENNAGATEAREA 0.0894 LAYER M8 ;
    ANTENNAGATEAREA 0.0894 LAYER M9 ;
    ANTENNAGATEAREA 0.0894 LAYER MRDL ;
  END CE1

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAGATEAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.142736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.142736 LAYER M2 ;
    ANTENNAMAXAREACAR 62.31165 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 69.52659 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 76.74104 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 83.95503 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[3]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.269224 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.269224 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.081 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56884 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56884 LAYER M2 ;
    ANTENNAMAXAREACAR 7.988725 LAYER M2 ;
    ANTENNAGATEAREA 0.081 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 9.859802 LAYER M3 ;
    ANTENNAGATEAREA 0.081 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 11.73076 LAYER M4 ;
    ANTENNAGATEAREA 0.081 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 13.60159 LAYER M5 ;
    ANTENNAGATEAREA 0.081 LAYER M6 ;
    ANTENNAGATEAREA 0.081 LAYER M7 ;
    ANTENNAGATEAREA 0.081 LAYER M8 ;
    ANTENNAGATEAREA 0.081 LAYER M9 ;
    ANTENNAGATEAREA 0.081 LAYER MRDL ;
  END OEB1

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.58662 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.58662 LAYER M2 ;
    ANTENNAMAXAREACAR 11.89816 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.93502 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.97181 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.00853 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.59904 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.59904 LAYER M2 ;
    ANTENNAMAXAREACAR 11.98317 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 13.02002 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.05681 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.09353 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.5160 52.1790 46.8160 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.6170 52.1790 9.9170 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.5160 52.1790 10.8170 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.1160 52.1790 23.4150 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.6140 52.1790 45.9150 52.4790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 69.7947 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 69.7947 LAYER M5 ;
  END VDDL

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.081 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56302 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56302 LAYER M2 ;
    ANTENNAMAXAREACAR 7.916873 LAYER M2 ;
    ANTENNAGATEAREA 0.081 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 9.787955 LAYER M3 ;
    ANTENNAGATEAREA 0.081 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 11.65891 LAYER M4 ;
    ANTENNAGATEAREA 0.081 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 13.52975 LAYER M5 ;
    ANTENNAGATEAREA 0.081 LAYER M6 ;
    ANTENNAGATEAREA 0.081 LAYER M7 ;
    ANTENNAGATEAREA 0.081 LAYER M8 ;
    ANTENNAGATEAREA 0.081 LAYER M9 ;
    ANTENNAGATEAREA 0.081 LAYER MRDL ;
  END OEB2

  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.9160 52.1790 7.2170 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.8170 52.1790 8.1170 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.8170 52.1790 17.1160 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.7170 52.1790 18.0170 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.3170 52.1790 48.6170 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.2170 52.1790 49.5160 52.4790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 92.8485 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 92.8485 LAYER M5 ;
  END VDD

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.295008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.295008 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.3262 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3262 LAYER M4 ;
    ANTENNAMAXAREACAR 15.01649 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 19.44825 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.43702 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43702 LAYER M4 ;
    ANTENNAMAXAREACAR 14.36045 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.50158 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.123568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.123568 LAYER M3 ;
    ANTENNAMAXAREACAR 33.06199 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.20189 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.34151 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.123568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.123568 LAYER M3 ;
    ANTENNAMAXAREACAR 33.06199 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.20189 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.34151 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 41.9970 55.6450 42.1970 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 41.9970 55.6450 42.1970 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 41.9970 55.6450 42.1970 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 41.9970 55.6450 42.1970 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 41.9970 55.6450 42.1970 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.2043 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.672754 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.672754 LAYER M2 ;
    ANTENNAMAXAREACAR 10.51521 LAYER M2 ;
    ANTENNAGATEAREA 0.6282 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.67607 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.67607 LAYER M3 ;
    ANTENNAMAXAREACAR 12.15055 LAYER M3 ;
    ANTENNAGATEAREA 0.6282 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 15.01542 LAYER M4 ;
    ANTENNAGATEAREA 0.6282 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.25576 LAYER M5 ;
    ANTENNAGATEAREA 0.6282 LAYER M6 ;
    ANTENNAGATEAREA 0.6282 LAYER M7 ;
    ANTENNAGATEAREA 0.6282 LAYER M8 ;
    ANTENNAGATEAREA 0.6282 LAYER M9 ;
    ANTENNAGATEAREA 0.6282 LAYER MRDL ;
  END SD

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 45.5510 55.6450 45.7510 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 45.5510 55.6450 45.7510 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 45.5510 55.6450 45.7510 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 45.5510 55.6450 45.7510 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 45.5510 55.6450 45.7510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.534885 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.534885 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 36.56684 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 39.6086 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.65017 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.5510 0.2000 45.7510 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 45.5510 0.2000 45.7510 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 45.5510 0.2000 45.7510 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 45.5510 0.2000 45.7510 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 45.5510 0.2000 45.7510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.587205 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.587205 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 37.99624 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 41.03791 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 44.07938 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 42.3370 55.6450 42.5370 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 42.3370 55.6450 42.5370 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 42.3370 55.6450 42.5370 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 42.3370 55.6450 42.5370 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 42.3370 55.6450 42.5370 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.54727 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.54727 LAYER M2 ;
    ANTENNAMAXAREACAR 27.62053 LAYER M2 ;
    ANTENNAGATEAREA 0.132 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.39759 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.39759 LAYER M3 ;
    ANTENNAMAXAREACAR 29.1118 LAYER M3 ;
    ANTENNAGATEAREA 0.132 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 46.92944 LAYER M4 ;
    ANTENNAGATEAREA 0.132 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 48.07483 LAYER M5 ;
    ANTENNAGATEAREA 0.132 LAYER M6 ;
    ANTENNAGATEAREA 0.132 LAYER M7 ;
    ANTENNAGATEAREA 0.132 LAYER M8 ;
    ANTENNAGATEAREA 0.132 LAYER M9 ;
    ANTENNAGATEAREA 0.132 LAYER MRDL ;
  END DS1

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 42.3370 0.2000 42.5370 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 42.3370 0.2000 42.5370 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 42.3370 0.2000 42.5370 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 42.3370 0.2000 42.5370 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 42.3370 0.2000 42.5370 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.5185 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5185 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.25657 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.25657 LAYER M2 ;
    ANTENNAMAXAREACAR 13.9726 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.154727 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.154727 LAYER M3 ;
    ANTENNAMAXAREACAR 27.75069 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 42.61741 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 45.93916 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS2

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28128 LAYER M3 ;
    ANTENNAMAXAREACAR 62.2616 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47654 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.691 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.270888 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.1660 52.1790 18.4670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.9670 52.1790 47.2660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.4660 52.1790 15.7660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.8660 52.1790 48.1660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.3660 52.1790 16.6670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.7660 52.1790 49.0670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.2660 52.1790 17.5670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.5670 52.1790 14.8660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.1670 52.1790 45.4670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.7670 52.1790 13.0670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.0660 52.1790 46.3660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.6660 52.1790 13.9660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.2660 52.1790 44.5660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8660 52.1790 12.1660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.3670 52.1790 43.6660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.5660 52.1790 32.8650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.9670 52.1790 11.2660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.4670 52.1790 42.7670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.6660 52.1790 31.9660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.0670 52.1790 10.3670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.5660 52.1790 41.8670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.7650 52.1790 31.0660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.1660 52.1790 9.4670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.8670 52.1790 39.1660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.0660 52.1790 28.3650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.4670 52.1790 6.7660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.9670 52.1790 38.2670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.1660 52.1790 27.4660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.5670 52.1790 5.8670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.7670 52.1790 40.0660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.9660 52.1790 29.2650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.3670 52.1790 7.6660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.6660 52.1790 40.9670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.8650 52.1790 30.1660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.2660 52.1790 8.5670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.2660 52.1790 35.5660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.4650 52.1790 24.7650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.8660 52.1790 3.1660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.3670 52.1790 34.6670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.5660 52.1790 23.8660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9670 52.1790 2.2670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.4660 52.1790 33.7660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.6650 52.1790 22.9650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.0650 52.1790 1.3650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.0660 52.1790 37.3670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.2650 52.1790 26.5660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.6660 52.1790 4.9670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.1660 52.1790 36.4670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.3650 52.1790 25.6660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.7660 52.1790 4.0670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.1650 52.1790 54.4650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.7650 52.1790 22.0650 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.3670 52.1790 52.6670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.9670 52.1790 20.2670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.2660 52.1790 53.5660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.8660 52.1790 21.1660 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.4670 52.1790 51.7670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.0670 52.1790 19.3670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.5660 52.1790 50.8670 52.4790 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.6660 52.1790 49.9670 52.4790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 24.258 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1662.414 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1662.414 LAYER M5 ;
    ANTENNAMAXAREACAR 159.2478 LAYER M5 ;
    ANTENNAGATEAREA 24.258 LAYER M6 ;
    ANTENNAGATEAREA 24.258 LAYER M7 ;
    ANTENNAGATEAREA 24.258 LAYER M8 ;
    ANTENNAGATEAREA 24.258 LAYER M9 ;
    ANTENNAGATEAREA 24.258 LAYER MRDL ;
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0000 43.1370 1.5010 44.9510 ;
      RECT 54.1440 43.1370 55.6450 44.9510 ;
      RECT 0.0000 30.6190 3.0010 30.6330 ;
      RECT 0.0000 36.4620 54.8450 39.4630 ;
      RECT 0.0000 40.8630 0.8000 41.7370 ;
      RECT 52.6440 33.5080 55.6450 33.5220 ;
      RECT 54.8450 40.8490 55.6450 41.3970 ;
      RECT 0.0000 32.0330 0.8000 32.1220 ;
      RECT 54.8450 32.0190 55.6450 32.1080 ;
      RECT 0.0000 18.0520 55.6450 25.3140 ;
      RECT 0.0000 46.3510 55.6450 52.4790 ;
      RECT 0.0000 18.0460 54.8450 25.3140 ;
      RECT 0.0000 18.0460 54.8450 25.3140 ;
      RECT 0.0000 18.0460 54.8450 25.3140 ;
      RECT 0.0000 18.0460 54.8450 18.0520 ;
      RECT 0.8000 16.1920 54.8450 18.0460 ;
      RECT 0.8000 16.1860 55.6450 16.1920 ;
      RECT 0.0000 0.0000 20.5070 9.1790 ;
      RECT 0.0000 0.0000 20.5070 0.8000 ;
      RECT 0.0000 10.5800 55.6450 16.1860 ;
      RECT 0.8000 10.5800 54.8450 18.0460 ;
      RECT 0.8000 10.5800 54.8450 18.0460 ;
      RECT 0.8000 10.5800 54.8450 18.0460 ;
      RECT 0.8000 10.5800 55.6450 16.1920 ;
      RECT 0.8000 10.5800 55.6450 16.1920 ;
      RECT 0.8000 10.5800 55.6450 16.1920 ;
      RECT 0.8000 10.5790 55.6450 16.1860 ;
      RECT 0.8000 10.5790 55.6450 10.5800 ;
      RECT 0.8000 9.1800 54.8450 10.5790 ;
      RECT 0.0000 25.3140 54.8450 25.3280 ;
      RECT 0.0000 18.0520 54.8450 25.3280 ;
      RECT 0.0000 18.0520 54.8450 25.3280 ;
      RECT 0.0000 18.0520 54.8450 25.3280 ;
      RECT 0.8000 25.3280 54.8450 26.7140 ;
      RECT 0.0000 9.1790 54.8450 9.1800 ;
      RECT 0.0000 0.8000 54.8450 9.1800 ;
      RECT 0.0000 0.8000 54.8450 9.1800 ;
      RECT 0.0000 0.8000 54.8450 9.1800 ;
      RECT 0.0000 0.8000 55.6450 9.1790 ;
      RECT 0.8000 0.8000 54.8450 10.5790 ;
      RECT 0.8000 0.8000 54.8450 10.5790 ;
      RECT 0.8000 0.8000 54.8450 10.5790 ;
      RECT 35.3390 0.0000 55.6450 9.1790 ;
      RECT 35.3390 0.0000 55.6450 0.8000 ;
      RECT 0.8000 41.7370 54.8450 46.3510 ;
      RECT 0.8000 41.7370 54.8450 46.3510 ;
      RECT 0.8000 41.7370 54.8450 46.3510 ;
      RECT 0.8000 41.7370 54.8450 46.3510 ;
      RECT 0.0000 26.7280 55.6450 30.6190 ;
      RECT 0.8000 32.0190 54.8450 32.0330 ;
      RECT 0.8000 26.7140 55.6450 30.6190 ;
      RECT 0.8000 26.7140 55.6450 30.6190 ;
      RECT 0.8000 26.7140 55.6450 30.6190 ;
      RECT 0.8000 25.3280 54.8450 30.6190 ;
      RECT 0.8000 25.3280 54.8450 30.6190 ;
      RECT 0.8000 25.3280 54.8450 30.6190 ;
      RECT 0.8000 26.7140 55.6450 26.7280 ;
      RECT 0.8000 39.4630 54.8450 52.4790 ;
      RECT 0.8000 40.8490 54.8450 46.3510 ;
      RECT 0.8000 40.8490 54.8450 46.3510 ;
      RECT 0.8000 40.8490 54.8450 46.3510 ;
      RECT 0.8000 39.4630 54.8450 46.3510 ;
      RECT 0.8000 40.8490 54.8450 44.9510 ;
      RECT 0.8000 40.8490 54.8450 44.9510 ;
      RECT 0.8000 40.8490 54.8450 44.9510 ;
      RECT 0.8000 40.8490 54.8450 44.9510 ;
      RECT 0.8000 39.4630 54.8450 44.9510 ;
      RECT 0.8000 39.4630 54.8450 44.9510 ;
      RECT 0.8000 39.4630 54.8450 44.9510 ;
      RECT 0.8000 39.4630 54.8450 44.9510 ;
      RECT 0.8000 39.4630 54.8450 43.1370 ;
      RECT 0.8000 41.3970 54.8450 41.7370 ;
      RECT 0.0000 33.5220 55.6450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6330 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 0.8000 30.6190 54.8450 39.4490 ;
      RECT 21.9070 0.0000 22.7950 0.8000 ;
    LAYER PO ;
      RECT 0.0000 0.0000 55.6450 52.4790 ;
    LAYER M4 ;
      RECT 0.9000 40.9490 54.7450 40.9630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 30.5330 54.7450 33.6080 ;
      RECT 0.9000 26.8140 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 0.0000 43.2370 1.5010 44.8510 ;
      RECT 0.0000 40.9630 0.9000 41.6370 ;
      RECT 54.1440 43.2370 55.6450 44.8510 ;
      RECT 54.7450 40.9490 55.6450 41.2970 ;
      RECT 0.0000 46.4510 55.6450 52.4790 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.0000 30.5190 54.7450 30.5330 ;
      RECT 0.0000 26.8280 54.7450 30.5330 ;
      RECT 0.0000 26.8280 55.6450 30.5190 ;
      RECT 0.0000 25.2140 54.7450 25.2280 ;
      RECT 0.0000 18.1460 54.7450 25.2280 ;
      RECT 0.0000 18.1460 54.7450 25.2280 ;
      RECT 0.0000 18.1520 55.6450 25.2140 ;
      RECT 0.0000 18.1460 54.7450 18.1520 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.0000 0.0000 20.4070 9.0800 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 44.8510 54.7450 46.4510 ;
      RECT 0.9000 43.2370 54.7450 44.8510 ;
      RECT 0.9000 41.6370 54.7450 43.2370 ;
      RECT 0.9000 41.2970 54.7450 41.6370 ;
      RECT 0.9000 40.9630 54.7450 41.2970 ;
    LAYER M3 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 0.0000 43.2370 1.5010 44.8510 ;
      RECT 0.0000 40.9630 0.9000 41.6370 ;
      RECT 54.1440 43.2370 55.6450 44.8510 ;
      RECT 54.7450 40.9490 55.6450 41.2970 ;
      RECT 0.0000 46.4510 55.6450 52.4790 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.0000 30.5190 54.7450 30.5330 ;
      RECT 0.0000 26.8280 54.7450 30.5330 ;
      RECT 0.0000 26.8280 55.6450 30.5190 ;
      RECT 0.0000 25.2140 54.7450 25.2280 ;
      RECT 0.0000 18.1460 54.7450 25.2280 ;
      RECT 0.0000 18.1460 54.7450 25.2280 ;
      RECT 0.0000 18.1520 55.6450 25.2140 ;
      RECT 0.0000 18.1460 54.7450 18.1520 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.0000 0.0000 20.4070 9.0800 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 44.8510 54.7450 46.4510 ;
      RECT 0.9000 43.2370 54.7450 44.8510 ;
      RECT 0.9000 41.6370 54.7450 43.2370 ;
      RECT 0.9000 41.2970 54.7450 41.6370 ;
      RECT 0.9000 40.9630 54.7450 41.2970 ;
      RECT 0.9000 40.9490 54.7450 40.9630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 30.5330 54.7450 33.6080 ;
      RECT 0.9000 26.8140 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
    LAYER M2 ;
      RECT 0.0000 40.9630 0.9000 41.6370 ;
      RECT 54.7450 40.9490 55.6450 41.2970 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 0.0000 43.2370 1.5010 44.8510 ;
      RECT 54.1440 43.2370 55.6450 44.8510 ;
      RECT 0.0000 46.4510 55.6450 52.4790 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.0000 30.5190 54.7450 30.5330 ;
      RECT 0.0000 26.8280 54.7450 30.5330 ;
      RECT 0.0000 26.8280 55.6450 30.5190 ;
      RECT 0.0000 25.2140 54.7450 25.2280 ;
      RECT 0.0000 18.1460 54.7450 25.2280 ;
      RECT 0.0000 18.1460 54.7450 25.2280 ;
      RECT 0.0000 18.1520 55.6450 25.2140 ;
      RECT 0.0000 18.1460 54.7450 18.1520 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.0000 0.0000 20.4070 9.0800 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 0.9000 54.7450 52.4790 ;
      RECT 0.9000 44.8510 54.7450 46.4510 ;
      RECT 0.9000 43.2370 54.7450 44.8510 ;
      RECT 0.9000 41.6370 54.7450 43.2370 ;
      RECT 0.9000 41.2970 54.7450 41.6370 ;
      RECT 0.9000 40.9630 54.7450 41.2970 ;
      RECT 0.9000 40.9490 54.7450 40.9630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 30.5330 54.7450 33.6080 ;
      RECT 0.9000 26.8140 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 16.0920 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 55.6450 52.4790 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 55.6450 52.4790 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 55.6450 52.4790 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 55.6450 52.4790 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 55.6450 52.4790 ;
    LAYER M5 ;
      RECT 0.0000 51.4790 0.3650 52.4790 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 55.1650 51.4790 55.6450 52.4790 ;
      RECT 0.0000 40.9630 0.9000 41.6370 ;
      RECT 0.0000 36.3620 54.7450 39.3630 ;
      RECT 0.0000 43.2370 1.5010 44.8510 ;
      RECT 54.1440 43.2370 55.6450 44.8510 ;
      RECT 54.7450 40.9490 55.6450 41.2970 ;
      RECT 0.0000 18.1520 55.6450 25.2140 ;
      RECT 0.9000 30.5330 54.7450 33.6080 ;
      RECT 0.0000 46.4510 55.6450 51.4790 ;
      RECT 0.9000 43.2370 54.7450 51.4790 ;
      RECT 0.9000 43.2370 54.7450 51.4790 ;
      RECT 0.9000 41.6370 54.7450 51.4790 ;
      RECT 0.0000 18.1460 54.7450 25.2140 ;
      RECT 0.0000 18.1460 54.7450 25.2140 ;
      RECT 0.0000 18.1460 54.7450 25.2140 ;
      RECT 0.0000 18.1460 54.7450 18.1520 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.0000 30.5190 54.7450 30.5330 ;
      RECT 0.0000 26.8280 54.7450 30.5330 ;
      RECT 0.0000 26.8280 55.6450 30.5190 ;
      RECT 0.0000 25.2140 54.7450 25.2280 ;
      RECT 0.0000 18.1520 54.7450 25.2280 ;
      RECT 0.0000 18.1520 54.7450 25.2280 ;
      RECT 0.0000 18.1520 54.7450 25.2280 ;
      RECT 0.9000 26.8280 54.7450 33.6080 ;
      RECT 0.9000 26.8140 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 30.5190 ;
      RECT 0.9000 25.2280 54.7450 30.5190 ;
      RECT 0.9000 25.2280 54.7450 30.5190 ;
      RECT 0.9000 25.2280 54.7450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.9000 10.6800 54.7450 18.1460 ;
      RECT 0.9000 10.6800 54.7450 18.1460 ;
      RECT 0.9000 10.6800 54.7450 18.1460 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.0000 0.0000 20.4070 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 30.5330 54.7450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 39.3630 54.7450 51.4790 ;
      RECT 0.9000 39.3630 54.7450 46.4510 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
      RECT 0.9000 39.3630 54.7450 43.2370 ;
  END
END SRAMLP2RW16x4

MACRO SRAMLP2RW16x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 65.407 BY 54.861 ;
  SYMMETRY X Y R90 ;

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.5450 0.0000 41.7450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.5450 0.0000 41.7450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.5450 0.0000 41.7450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.5450 0.0000 41.7450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.5450 0.0000 41.7450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[2]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.9130 0.0000 43.1130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.9130 0.0000 43.1130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.9130 0.0000 43.1130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.9130 0.0000 43.1130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.9130 0.0000 43.1130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[3]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0800 0.0000 44.2800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0800 0.0000 44.2800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0800 0.0000 44.2800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0800 0.0000 44.2800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0800 0.0000 44.2800 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[5]

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 44.5960 65.4070 44.7960 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 44.5960 65.4070 44.7960 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 44.5960 65.4070 44.7960 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 44.5960 65.4070 44.7960 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 44.5960 65.4070 44.7960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
  END DS1

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    ANTENNADIFFAREA 1.84416 LAYER M3 ;
    ANTENNADIFFAREA 1.84416 LAYER M4 ;
    ANTENNADIFFAREA 1.84416 LAYER M5 ;
    ANTENNADIFFAREA 1.84416 LAYER M6 ;
    ANTENNADIFFAREA 1.84416 LAYER M7 ;
    ANTENNADIFFAREA 1.84416 LAYER M8 ;
    ANTENNADIFFAREA 1.84416 LAYER M9 ;
    ANTENNADIFFAREA 1.84416 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.1716 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.07152 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.07152 LAYER M3 ;
    ANTENNAMAXAREACAR 24.99403 LAYER M3 ;
    ANTENNAGATEAREA 0.1716 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M4 ;
    ANTENNAMAXAREACAR 32.06142 LAYER M4 ;
    ANTENNAGATEAREA 0.1716 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M5 ;
    ANTENNAMAXAREACAR 39.12876 LAYER M5 ;
    ANTENNAGATEAREA 0.1716 LAYER M6 ;
    ANTENNAGATEAREA 0.1716 LAYER M7 ;
    ANTENNAGATEAREA 0.1716 LAYER M8 ;
    ANTENNAGATEAREA 0.1716 LAYER M9 ;
    ANTENNAGATEAREA 0.1716 LAYER MRDL ;
  END O2[0]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 9.8030 65.4070 10.0030 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 9.8030 65.4070 10.0030 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 9.8030 65.4070 10.0030 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 9.8030 65.4070 10.0030 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 9.8030 65.4070 10.0030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15418 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15418 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.558163 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.558163 LAYER M2 ;
    ANTENNAMAXAREACAR 11.70338 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.74025 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.77706 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.8138 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8040 0.2000 10.0040 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8040 0.2000 10.0040 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8040 0.2000 10.0040 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8040 0.2000 10.0040 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8040 0.2000 10.0040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15418 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15418 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.55662 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.55662 LAYER M2 ;
    ANTENNAMAXAREACAR 11.69282 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.72969 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.7665 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.80324 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 44.2560 65.4070 44.4560 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 44.2560 65.4070 44.4560 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 44.2560 65.4070 44.4560 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 44.2560 65.4070 44.4560 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 44.2560 65.4070 44.4560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.2256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.804608 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.804608 LAYER M2 ;
    ANTENNAMAXAREACAR 8.542707 LAYER M2 ;
    ANTENNAGATEAREA 0.2256 LAYER M3 ;
    ANTENNAGATEAREA 0.2256 LAYER M4 ;
    ANTENNAGATEAREA 0.2256 LAYER M5 ;
    ANTENNAGATEAREA 0.2256 LAYER M6 ;
    ANTENNAGATEAREA 0.2256 LAYER M7 ;
    ANTENNAGATEAREA 0.2256 LAYER M8 ;
    ANTENNAGATEAREA 0.2256 LAYER M9 ;
    ANTENNAGATEAREA 0.2256 LAYER MRDL ;
  END SD

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 47.8100 65.4070 48.0100 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 47.8100 65.4070 48.0100 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 47.8100 65.4070 48.0100 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 47.8100 65.4070 48.0100 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 47.8100 65.4070 48.0100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.324765 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.324765 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 30.82629 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 33.86844 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.91038 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 44.6120 0.2000 44.8120 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 44.6120 0.2000 44.8120 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 44.6120 0.2000 44.8120 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 44.6120 0.2000 44.8120 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 44.6120 0.2000 44.8120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.34288 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.34288 LAYER M1 ;
    ANTENNAGATEAREA 0.2256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.443613 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.443613 LAYER M2 ;
    ANTENNAMAXAREACAR 6.902549 LAYER M2 ;
    ANTENNAGATEAREA 0.8058 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 8.112283 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.112283 LAYER M3 ;
    ANTENNAMAXAREACAR 46.67783 LAYER M3 ;
    ANTENNAGATEAREA 0.8058 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 18.3684 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3684 LAYER M4 ;
    ANTENNAMAXAREACAR 69.47304 LAYER M4 ;
    ANTENNAGATEAREA 0.8058 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 97.5558 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 97.5558 LAYER M5 ;
    ANTENNAMAXAREACAR 190.54 LAYER M5 ;
    ANTENNAGATEAREA 0.8058 LAYER M6 ;
    ANTENNAGATEAREA 0.8058 LAYER M7 ;
    ANTENNAGATEAREA 0.8058 LAYER M8 ;
    ANTENNAGATEAREA 0.8058 LAYER M9 ;
    ANTENNAGATEAREA 0.8058 LAYER MRDL ;
  END DS2

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 47.8260 0.2000 48.0260 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 47.8260 0.2000 48.0260 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 47.8260 0.2000 48.0260 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 47.8260 0.2000 48.0260 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 47.8260 0.2000 48.0260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.437625 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.437625 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 33.90966 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.95161 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 39.99334 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.3990 0.0000 20.5990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.3990 0.0000 20.5990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.3990 0.0000 20.5990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.3990 0.0000 20.5990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.3990 0.0000 20.5990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.897997 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.897997 LAYER M2 ;
    ANTENNAMAXAREACAR 7.228198 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.284904 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.341539 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.39811 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7750 0.0000 44.9750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7750 0.0000 44.9750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7750 0.0000 44.9750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7750 0.0000 44.9750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7750 0.0000 44.9750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.903817 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.903817 LAYER M2 ;
    ANTENNAMAXAREACAR 7.268784 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.325487 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.38212 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.43868 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB1

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.1990 0.0000 30.3990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.1990 0.0000 30.3990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.1990 0.0000 30.3990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.1990 0.0000 30.3990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.1990 0.0000 30.3990 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[2]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.4020 0.0000 35.6020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.4020 0.0000 35.6020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.4020 0.0000 35.6020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.4020 0.0000 35.6020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.4020 0.0000 35.6020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[7]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.7700 0.0000 36.9700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.7700 0.0000 36.9700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.7700 0.0000 36.9700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.7700 0.0000 36.9700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.7700 0.0000 36.9700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[1]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.1380 0.0000 38.3380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.1380 0.0000 38.3380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.1380 0.0000 38.3380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.1380 0.0000 38.3380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.1380 0.0000 38.3380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[6]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.5060 0.0000 39.7060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.5060 0.0000 39.7060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.5060 0.0000 39.7060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.5060 0.0000 39.7060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.5060 0.0000 39.7060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[4]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.8740 0.0000 41.0740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.8740 0.0000 41.0740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.8740 0.0000 41.0740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.8740 0.0000 41.0740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.8740 0.0000 41.0740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.2420 0.0000 42.4420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.2420 0.0000 42.4420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.2420 0.0000 42.4420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.2420 0.0000 42.4420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.2420 0.0000 42.4420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[3]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.6100 0.0000 43.8100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.6100 0.0000 43.8100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.6100 0.0000 43.8100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.6100 0.0000 43.8100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.6100 0.0000 43.8100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I1[5]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.7270 0.0000 24.9270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.7270 0.0000 24.9270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.7270 0.0000 24.9270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.7270 0.0000 24.9270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.7270 0.0000 24.9270 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[7]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[1]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.4630 0.0000 27.6630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.4630 0.0000 27.6630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.4630 0.0000 27.6630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.4630 0.0000 27.6630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.4630 0.0000 27.6630 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[6]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.8310 0.0000 29.0310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.8310 0.0000 29.0310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.8310 0.0000 29.0310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.8310 0.0000 29.0310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.8310 0.0000 29.0310 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[4]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.5670 0.0000 31.7670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.5670 0.0000 31.7670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.5670 0.0000 31.7670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.5670 0.0000 31.7670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.5670 0.0000 31.7670 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[3]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[5]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.7050 0.0000 34.9050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.7050 0.0000 34.9050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.7050 0.0000 34.9050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.7050 0.0000 34.9050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.7050 0.0000 34.9050 0.2000 ;
    END
    ANTENNADIFFAREA 1.9074 LAYER M3 ;
    ANTENNADIFFAREA 1.9074 LAYER M4 ;
    ANTENNADIFFAREA 1.9074 LAYER M5 ;
    ANTENNADIFFAREA 1.9074 LAYER M6 ;
    ANTENNADIFFAREA 1.9074 LAYER M7 ;
    ANTENNADIFFAREA 1.9074 LAYER M8 ;
    ANTENNADIFFAREA 1.9074 LAYER M9 ;
    ANTENNADIFFAREA 1.9074 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.2844 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.06294 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.06294 LAYER M3 ;
    ANTENNAMAXAREACAR 21.91653 LAYER M3 ;
    ANTENNAGATEAREA 0.2844 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M4 ;
    ANTENNAMAXAREACAR 26.18076 LAYER M4 ;
    ANTENNAGATEAREA 0.2844 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M5 ;
    ANTENNAMAXAREACAR 30.44497 LAYER M5 ;
    ANTENNAGATEAREA 0.2844 LAYER M6 ;
    ANTENNAGATEAREA 0.2844 LAYER M7 ;
    ANTENNAGATEAREA 0.2844 LAYER M8 ;
    ANTENNAGATEAREA 0.2844 LAYER M9 ;
    ANTENNAGATEAREA 0.2844 LAYER MRDL ;
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.0730 0.0000 36.2730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.0730 0.0000 36.2730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.0730 0.0000 36.2730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.0730 0.0000 36.2730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.0730 0.0000 36.2730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[7]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.4410 0.0000 37.6410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.4410 0.0000 37.6410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.4410 0.0000 37.6410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.4410 0.0000 37.6410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.4410 0.0000 37.6410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[1]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.8090 0.0000 39.0090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.8090 0.0000 39.0090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.8090 0.0000 39.0090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.8090 0.0000 39.0090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.8090 0.0000 39.0090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[6]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.1770 0.0000 40.3770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.1770 0.0000 40.3770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.1770 0.0000 40.3770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.1770 0.0000 40.3770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.1770 0.0000 40.3770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[4]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.2760 0.2000 17.4760 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.2760 0.2000 17.4760 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.2760 0.2000 17.4760 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.2760 0.2000 17.4760 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.2760 0.2000 17.4760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.1128 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.65322 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.65322 LAYER M4 ;
    ANTENNAMAXAREACAR 22.67857 LAYER M4 ;
    ANTENNAGATEAREA 28.8444 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 2044.503 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2044.503 LAYER M5 ;
    ANTENNAMAXAREACAR 186.1565 LAYER M5 ;
    ANTENNAGATEAREA 28.8444 LAYER M6 ;
    ANTENNAGATEAREA 28.8444 LAYER M7 ;
    ANTENNAGATEAREA 28.8444 LAYER M8 ;
    ANTENNAGATEAREA 28.8444 LAYER M9 ;
    ANTENNAGATEAREA 28.8444 LAYER MRDL ;
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8160 0.2000 17.0160 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8160 0.2000 17.0160 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8160 0.2000 17.0160 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8160 0.2000 17.0160 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8160 0.2000 17.0160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.39514 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.39514 LAYER M4 ;
    ANTENNAMAXAREACAR 13.94555 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.0867 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 17.2760 65.4070 17.4760 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 17.2760 65.4070 17.4760 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 17.2760 65.4070 17.4760 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 17.2760 65.4070 17.4760 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 17.2760 65.4070 17.4760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.1128 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.70704 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.70704 LAYER M4 ;
    ANTENNAMAXAREACAR 22.97495 LAYER M4 ;
    ANTENNAGATEAREA 0.1128 LAYER M5 ;
    ANTENNAGATEAREA 0.1128 LAYER M6 ;
    ANTENNAGATEAREA 0.1128 LAYER M7 ;
    ANTENNAGATEAREA 0.1128 LAYER M8 ;
    ANTENNAGATEAREA 0.1128 LAYER M9 ;
    ANTENNAGATEAREA 0.1128 LAYER MRDL ;
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 16.8160 65.4070 17.0160 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 16.8160 65.4070 17.0160 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 16.8160 65.4070 17.0160 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 16.8160 65.4070 17.0160 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 16.8160 65.4070 17.0160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.39652 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.39652 LAYER M4 ;
    ANTENNAMAXAREACAR 13.98325 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.12441 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 42.2560 65.4070 42.4560 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 42.2560 65.4070 42.4560 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 42.2560 65.4070 42.4560 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 42.2560 65.4070 42.4560 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 42.2560 65.4070 42.4560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 34.9150 65.4070 35.1150 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 34.9150 65.4070 35.1150 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 34.9150 65.4070 35.1150 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 34.9150 65.4070 35.1150 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 34.9150 65.4070 35.1150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 33.4260 65.4070 33.6260 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 33.4260 65.4070 33.6260 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 33.4260 65.4070 33.6260 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 33.4260 65.4070 33.6260 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 33.4260 65.4070 33.6260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2070 28.1210 65.4070 28.3210 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2070 28.1210 65.4070 28.3210 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2070 28.1210 65.4070 28.3210 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2070 28.1210 65.4070 28.3210 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2070 28.1210 65.4070 28.3210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAGATEAREA 0.2748 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 4.348947 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.348947 LAYER M2 ;
    ANTENNAMAXAREACAR 27.14591 LAYER M2 ;
    ANTENNAGATEAREA 0.2748 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.69579 LAYER M3 ;
    ANTENNAGATEAREA 0.2748 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 28.24564 LAYER M4 ;
    ANTENNAGATEAREA 0.2748 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 28.79545 LAYER M5 ;
    ANTENNAGATEAREA 0.2748 LAYER M6 ;
    ANTENNAGATEAREA 0.2748 LAYER M7 ;
    ANTENNAGATEAREA 0.2748 LAYER M8 ;
    ANTENNAGATEAREA 0.2748 LAYER M9 ;
    ANTENNAGATEAREA 0.2748 LAYER MRDL ;
  END A1[3]

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 57.5280 54.5610 57.8270 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.4290 54.5610 58.7280 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.8280 54.5610 19.1290 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.0290 54.5610 8.3290 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.1280 54.5610 7.4290 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.7290 54.5610 20.0290 54.8610 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 97.1022 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 97.1022 LAYER M5 ;
  END VDDL

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.168 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 10.52672 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.52672 LAYER M3 ;
    ANTENNAMAXAREACAR 63.90732 LAYER M3 ;
    ANTENNAGATEAREA 0.5532 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 14.45952 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.45952 LAYER M4 ;
    ANTENNAMAXAREACAR 39.38992 LAYER M4 ;
    ANTENNAGATEAREA 0.5532 LAYER M5 ;
    ANTENNAGATEAREA 0.5532 LAYER M6 ;
    ANTENNAGATEAREA 0.5532 LAYER M7 ;
    ANTENNAGATEAREA 0.5532 LAYER M8 ;
    ANTENNAGATEAREA 0.5532 LAYER M9 ;
    ANTENNAGATEAREA 0.5532 LAYER MRDL ;
  END I2[0]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[7]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[1]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[6]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.1600 0.0000 28.3600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.1600 0.0000 28.3600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.1600 0.0000 28.3600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.1600 0.0000 28.3600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.1600 0.0000 28.3600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[4]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.5280 0.0000 29.7280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.5280 0.0000 29.7280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.5280 0.0000 29.7280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.5280 0.0000 29.7280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.5280 0.0000 29.7280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.8960 0.0000 31.0960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.8960 0.0000 31.0960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.8960 0.0000 31.0960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.8960 0.0000 31.0960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.8960 0.0000 31.0960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[3]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.2640 0.0000 32.4640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.2640 0.0000 32.4640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.2640 0.0000 32.4640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.2640 0.0000 32.4640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.2640 0.0000 32.4640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END I2[5]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.0340 0.0000 34.2340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.0340 0.0000 34.2340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.0340 0.0000 34.2340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.0340 0.0000 34.2340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.0340 0.0000 34.2340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.168 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 10.52672 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.52672 LAYER M3 ;
    ANTENNAMAXAREACAR 63.90732 LAYER M3 ;
    ANTENNAGATEAREA 0.5532 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 14.17725 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.17725 LAYER M4 ;
    ANTENNAMAXAREACAR 38.87968 LAYER M4 ;
    ANTENNAGATEAREA 0.5532 LAYER M5 ;
    ANTENNAGATEAREA 0.5532 LAYER M6 ;
    ANTENNAGATEAREA 0.5532 LAYER M7 ;
    ANTENNAGATEAREA 0.5532 LAYER M8 ;
    ANTENNAGATEAREA 0.5532 LAYER M9 ;
    ANTENNAGATEAREA 0.5532 LAYER MRDL ;
  END I1[0]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.1210 0.2000 28.3210 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 28.1210 0.2000 28.3210 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 28.1210 0.2000 28.3210 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 28.1210 0.2000 28.3210 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 28.1210 0.2000 28.3210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAGATEAREA 0.2748 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 4.32806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.32806 LAYER M2 ;
    ANTENNAMAXAREACAR 27.1349 LAYER M2 ;
    ANTENNAGATEAREA 0.2748 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.68478 LAYER M3 ;
    ANTENNAGATEAREA 0.2748 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 28.23463 LAYER M4 ;
    ANTENNAGATEAREA 0.2748 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 28.78444 LAYER M5 ;
    ANTENNAGATEAREA 0.2748 LAYER M6 ;
    ANTENNAGATEAREA 0.2748 LAYER M7 ;
    ANTENNAGATEAREA 0.2748 LAYER M8 ;
    ANTENNAGATEAREA 0.2748 LAYER M9 ;
    ANTENNAGATEAREA 0.2748 LAYER MRDL ;
  END A2[3]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 42.2560 0.2000 42.4560 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 42.2560 0.2000 42.4560 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 42.2560 0.2000 42.4560 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 42.2560 0.2000 42.4560 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 42.2560 0.2000 42.4560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 34.9150 0.2000 35.1150 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 34.9150 0.2000 35.1150 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 34.9150 0.2000 35.1150 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 34.9150 0.2000 35.1150 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 34.9150 0.2000 35.1150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 33.4260 0.2000 33.6260 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 33.4260 0.2000 33.6260 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 33.4260 0.2000 33.6260 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 33.4260 0.2000 33.6260 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 33.4260 0.2000 33.6260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 19.59 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 26.00353 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.00353 LAYER M3 ;
    ANTENNAMAXAREACAR 16.81964 LAYER M3 ;
    ANTENNAGATEAREA 19.59 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 72.7251 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 72.7251 LAYER M4 ;
    ANTENNAMAXAREACAR 20.53199 LAYER M4 ;
    ANTENNAGATEAREA 19.59 LAYER M5 ;
    ANTENNAGATEAREA 19.59 LAYER M6 ;
    ANTENNAGATEAREA 19.59 LAYER M7 ;
    ANTENNAGATEAREA 19.59 LAYER M8 ;
    ANTENNAGATEAREA 19.59 LAYER M9 ;
    ANTENNAGATEAREA 19.59 LAYER MRDL ;
  END A2[2]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 61.1280 54.5610 61.4270 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.0280 54.5610 62.3270 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.3280 54.5610 14.6280 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.2280 54.5610 15.5280 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.1290 54.5610 16.4290 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.3290 54.5610 5.6280 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.4290 54.5610 4.7280 54.8610 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 2.1790 54.5610 2.4790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.6790 54.5610 6.9780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.5790 54.5610 7.8780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.2790 54.5610 10.5790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.1790 54.5610 11.4780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.4780 54.5610 8.7790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.3780 54.5610 9.6790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.7790 54.5610 6.0790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.3780 54.5610 18.6790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.4780 54.5610 17.7790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.5780 54.5610 16.8790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.6780 54.5610 15.9780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.7790 54.5610 15.0780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.8780 54.5610 14.1780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.9790 54.5610 13.2790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.0780 54.5610 12.3780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.6780 54.5610 24.9790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.9780 54.5610 22.2790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.7790 54.5610 24.0780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.8790 54.5610 23.1790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.2790 54.5610 19.5790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.3780 54.5610 36.6790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.1780 54.5610 38.4780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.1780 54.5610 47.4780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.9780 54.5610 49.2770 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.0790 54.5610 48.3790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.5790 54.5610 34.8780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.6780 54.5610 42.9780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.2780 54.5610 46.5780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.8790 54.5610 50.1800 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.0790 54.5610 39.3790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.5790 54.5610 43.8790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.3790 54.5610 45.6800 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.4780 54.5610 44.7770 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.9780 54.5610 40.2770 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.7780 54.5610 42.0780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.8790 54.5610 41.1800 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.0790 54.5610 30.3780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.8780 54.5610 32.1790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.3780 54.5610 63.6780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.7790 54.5610 60.0790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.1790 54.5610 56.4790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.5790 54.5610 52.8790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.7780 54.5610 51.0780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.2770 54.5610 64.5770 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.4770 54.5610 62.7770 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.5780 54.5610 61.8780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.6780 54.5610 60.9780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.8780 54.5610 59.1780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.9780 54.5610 58.2780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.0780 54.5610 57.3780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.2780 54.5610 55.5780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.3780 54.5610 54.6780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.4780 54.5610 53.7780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.6780 54.5610 51.9780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.6790 54.5610 33.9780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.7790 54.5610 33.0790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.5780 54.5610 25.8780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.9780 54.5610 31.2790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.4790 54.5610 26.7790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.2780 54.5610 37.5780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.4780 54.5610 35.7790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.3780 54.5610 27.6780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.2790 54.5610 28.5790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.1790 54.5610 29.4780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.0780 54.5610 21.3780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.1790 54.5610 20.4790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.8780 54.5610 5.1790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.9780 54.5610 4.2790 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.0780 54.5610 3.3780 54.8610 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.2780 54.5610 1.5780 54.8610 ;
    END
  END VSS
  OBS
    LAYER M3 ;
      RECT 0.9000 48.7100 65.4070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 48.7100 65.4070 48.7260 ;
      RECT 0.9000 47.1260 64.5070 48.7100 ;
      RECT 21.2990 0.0000 21.9880 0.9000 ;
      RECT 0.0000 45.5120 1.5010 47.1260 ;
      RECT 0.0000 43.1560 0.9000 43.9120 ;
      RECT 63.9060 45.4960 65.4070 47.1100 ;
      RECT 64.5070 43.1560 65.4070 43.5560 ;
      RECT 0.0000 35.8150 65.4070 41.5560 ;
      RECT 0.0000 29.0210 65.4070 32.7260 ;
      RECT 0.0000 18.1760 65.4070 27.4210 ;
      RECT 0.0000 10.7040 65.4070 16.1160 ;
      RECT 0.0000 0.0000 19.6990 9.1040 ;
      RECT 0.0000 9.1030 64.5070 9.1040 ;
      RECT 0.0000 0.9000 64.5070 9.1040 ;
      RECT 0.0000 0.9000 65.4070 9.1030 ;
      RECT 0.0000 0.0000 19.6990 0.9000 ;
      RECT 0.9000 47.1100 64.5070 47.1260 ;
      RECT 0.9000 45.5120 64.5070 47.1100 ;
      RECT 0.9000 45.4960 64.5070 45.5120 ;
      RECT 0.9000 43.9120 64.5070 45.4960 ;
      RECT 0.9000 43.5560 64.5070 43.9120 ;
      RECT 0.9000 43.1560 64.5070 43.5560 ;
      RECT 0.9000 41.5560 64.5070 43.1560 ;
      RECT 0.9000 32.7260 64.5070 35.8150 ;
      RECT 0.9000 27.4210 64.5070 29.0210 ;
      RECT 0.9000 16.1160 64.5070 18.1760 ;
      RECT 0.9000 10.7030 65.4070 16.1160 ;
      RECT 0.9000 10.7030 65.4070 10.7040 ;
      RECT 0.9000 9.1040 64.5070 10.7030 ;
      RECT 45.6750 0.0000 65.4070 9.1030 ;
      RECT 45.6750 0.0000 65.4070 0.9000 ;
      RECT 0.0000 48.7260 65.4070 54.8610 ;
    LAYER M2 ;
      RECT 0.0000 43.1560 0.9000 43.9120 ;
      RECT 64.5070 43.1560 65.4070 43.5560 ;
      RECT 21.2990 0.0000 21.9880 0.9000 ;
      RECT 0.0000 45.5120 1.5010 47.1260 ;
      RECT 63.9060 45.4960 65.4070 47.1100 ;
      RECT 0.0000 35.8150 65.4070 41.5560 ;
      RECT 0.0000 29.0210 65.4070 32.7260 ;
      RECT 0.0000 18.1760 65.4070 27.4210 ;
      RECT 0.0000 10.7040 65.4070 16.1160 ;
      RECT 0.0000 0.0000 19.6990 9.1040 ;
      RECT 0.0000 9.1030 64.5070 9.1040 ;
      RECT 0.0000 0.9000 64.5070 9.1040 ;
      RECT 0.0000 0.9000 65.4070 9.1030 ;
      RECT 0.0000 0.0000 19.6990 0.9000 ;
      RECT 0.9000 47.1100 64.5070 47.1260 ;
      RECT 0.9000 45.5120 64.5070 47.1100 ;
      RECT 0.9000 45.4960 64.5070 45.5120 ;
      RECT 0.9000 43.9120 64.5070 45.4960 ;
      RECT 0.9000 43.5560 64.5070 43.9120 ;
      RECT 0.9000 43.1560 64.5070 43.5560 ;
      RECT 0.9000 41.5560 64.5070 43.1560 ;
      RECT 0.9000 32.7260 64.5070 35.8150 ;
      RECT 0.9000 27.4210 64.5070 29.0210 ;
      RECT 0.9000 16.1160 64.5070 18.1760 ;
      RECT 0.9000 10.7030 65.4070 16.1160 ;
      RECT 0.9000 10.7030 65.4070 10.7040 ;
      RECT 0.9000 9.1040 64.5070 10.7030 ;
      RECT 45.6750 0.0000 65.4070 9.1030 ;
      RECT 45.6750 0.0000 65.4070 0.9000 ;
      RECT 0.0000 48.7260 65.4070 54.8610 ;
      RECT 0.9000 48.7100 65.4070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 48.7100 65.4070 48.7260 ;
      RECT 0.9000 47.1260 64.5070 48.7100 ;
    LAYER M1 ;
      RECT 0.0000 34.2260 0.8000 34.3150 ;
      RECT 64.6070 34.2260 65.4070 34.3150 ;
      RECT 0.0000 43.0560 0.8000 44.0120 ;
      RECT 64.6070 43.0560 65.4070 43.6560 ;
      RECT 21.1990 0.0000 22.0880 0.8000 ;
      RECT 0.0000 45.4120 1.5010 47.2260 ;
      RECT 63.9060 45.3960 65.4070 47.2100 ;
      RECT 0.0000 35.7150 65.4070 41.6560 ;
      RECT 0.0000 28.9210 65.4070 32.8260 ;
      RECT 0.0000 18.0760 65.4070 27.5210 ;
      RECT 0.0000 10.6040 65.4070 16.2160 ;
      RECT 0.0000 0.0000 19.7990 9.2040 ;
      RECT 0.0000 9.2030 64.6070 9.2040 ;
      RECT 0.0000 0.8000 64.6070 9.2040 ;
      RECT 0.0000 0.8000 65.4070 9.2030 ;
      RECT 0.0000 0.0000 19.7990 0.8000 ;
      RECT 0.8000 47.2100 64.6070 47.2260 ;
      RECT 0.8000 45.4120 64.6070 47.2100 ;
      RECT 0.8000 45.3960 64.6070 45.4120 ;
      RECT 0.8000 44.0120 64.6070 45.3960 ;
      RECT 0.8000 43.6560 64.6070 44.0120 ;
      RECT 0.8000 43.0560 64.6070 43.6560 ;
      RECT 0.8000 41.6560 64.6070 43.0560 ;
      RECT 0.8000 34.3150 64.6070 35.7150 ;
      RECT 0.8000 34.2260 64.6070 34.3150 ;
      RECT 0.8000 32.8260 64.6070 34.2260 ;
      RECT 0.8000 27.5210 64.6070 28.9210 ;
      RECT 0.8000 16.2160 64.6070 18.0760 ;
      RECT 0.8000 10.6030 65.4070 16.2160 ;
      RECT 0.8000 10.6030 65.4070 10.6040 ;
      RECT 0.8000 9.2040 64.6070 10.6030 ;
      RECT 45.5750 0.0000 65.4070 9.2030 ;
      RECT 45.5750 0.0000 65.4070 0.8000 ;
      RECT 0.0000 48.6260 65.4070 54.8610 ;
      RECT 0.8000 48.6100 65.4070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 0.8000 64.6070 54.8610 ;
      RECT 0.8000 48.6100 65.4070 48.6260 ;
      RECT 0.8000 47.2260 64.6070 48.6100 ;
    LAYER PO ;
      RECT 0.0000 0.0000 65.4070 54.8610 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 65.4070 54.8610 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 65.4070 54.8610 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 65.4070 54.8610 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 65.4070 54.8610 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 65.4070 54.8610 ;
    LAYER M5 ;
      RECT 65.2770 53.8610 65.4070 54.8610 ;
      RECT 0.0000 53.8610 0.5780 54.8610 ;
      RECT 21.2990 0.0000 21.9880 0.9000 ;
      RECT 0.0000 45.5120 1.5010 47.1260 ;
      RECT 0.0000 43.1560 0.9000 43.9120 ;
      RECT 63.9060 45.4960 65.4070 47.1100 ;
      RECT 64.5070 43.1560 65.4070 43.5560 ;
      RECT 0.0000 35.8150 65.4070 41.5560 ;
      RECT 0.0000 29.0210 65.4070 32.7260 ;
      RECT 0.0000 18.1760 65.4070 27.4210 ;
      RECT 0.0000 10.7040 65.4070 16.1160 ;
      RECT 0.0000 0.0000 19.6990 9.1040 ;
      RECT 0.0000 9.1030 64.5070 9.1040 ;
      RECT 0.0000 0.9000 64.5070 9.1040 ;
      RECT 0.0000 0.9000 65.4070 9.1030 ;
      RECT 0.0000 0.0000 19.6990 0.9000 ;
      RECT 0.9000 47.1100 64.5070 47.1260 ;
      RECT 0.9000 45.5120 64.5070 47.1100 ;
      RECT 0.9000 45.4960 64.5070 45.5120 ;
      RECT 0.9000 43.9120 64.5070 45.4960 ;
      RECT 0.9000 43.5560 64.5070 43.9120 ;
      RECT 0.9000 43.1560 64.5070 43.5560 ;
      RECT 0.9000 41.5560 64.5070 43.1560 ;
      RECT 0.9000 32.7260 64.5070 35.8150 ;
      RECT 0.9000 27.4210 64.5070 29.0210 ;
      RECT 0.9000 16.1160 64.5070 18.1760 ;
      RECT 0.9000 10.7030 65.4070 16.1160 ;
      RECT 0.9000 10.7030 65.4070 10.7040 ;
      RECT 0.9000 9.1040 64.5070 10.7030 ;
      RECT 45.6750 0.0000 65.4070 9.1030 ;
      RECT 45.6750 0.0000 65.4070 0.9000 ;
      RECT 0.0000 48.7260 65.4070 53.8610 ;
      RECT 0.9000 48.7100 65.4070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 0.9000 64.5070 53.8610 ;
      RECT 0.9000 48.7100 65.4070 48.7260 ;
      RECT 0.9000 47.1260 64.5070 48.7100 ;
    LAYER M4 ;
      RECT 21.2990 0.0000 21.9880 0.9000 ;
      RECT 0.0000 45.5120 1.5010 47.1260 ;
      RECT 0.0000 43.1560 0.9000 43.9120 ;
      RECT 63.9060 45.4960 65.4070 47.1100 ;
      RECT 64.5070 43.1560 65.4070 43.5560 ;
      RECT 0.0000 35.8150 65.4070 41.5560 ;
      RECT 0.0000 29.0210 65.4070 32.7260 ;
      RECT 0.0000 18.1760 65.4070 27.4210 ;
      RECT 0.0000 10.7040 65.4070 16.1160 ;
      RECT 0.0000 0.0000 19.6990 9.1040 ;
      RECT 0.0000 9.1030 64.5070 9.1040 ;
      RECT 0.0000 0.9000 64.5070 9.1040 ;
      RECT 0.0000 0.9000 65.4070 9.1030 ;
      RECT 0.0000 0.0000 19.6990 0.9000 ;
      RECT 0.9000 47.1100 64.5070 47.1260 ;
      RECT 0.9000 45.5120 64.5070 47.1100 ;
      RECT 0.9000 45.4960 64.5070 45.5120 ;
      RECT 0.9000 43.9120 64.5070 45.4960 ;
      RECT 0.9000 43.5560 64.5070 43.9120 ;
      RECT 0.9000 43.1560 64.5070 43.5560 ;
      RECT 0.9000 41.5560 64.5070 43.1560 ;
      RECT 0.9000 32.7260 64.5070 35.8150 ;
      RECT 0.9000 27.4210 64.5070 29.0210 ;
      RECT 0.9000 16.1160 64.5070 18.1760 ;
      RECT 0.9000 10.7030 65.4070 16.1160 ;
      RECT 0.9000 10.7030 65.4070 10.7040 ;
      RECT 0.9000 9.1040 64.5070 10.7030 ;
      RECT 45.6750 0.0000 65.4070 9.1030 ;
      RECT 45.6750 0.0000 65.4070 0.9000 ;
      RECT 0.0000 48.7260 65.4070 54.8610 ;
      RECT 0.9000 48.7100 65.4070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 0.9000 64.5070 54.8610 ;
      RECT 0.9000 48.7100 65.4070 48.7260 ;
      RECT 0.9000 47.1260 64.5070 48.7100 ;
  END
END SRAMLP2RW16x8

MACRO SRAMLP2RW16x16
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 87.653 BY 59.155 ;
  SYMMETRY X Y R90 ;

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 46.5730 0.2000 46.7730 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 46.5730 0.2000 46.7730 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 46.5730 0.2000 46.7730 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 46.5730 0.2000 46.7730 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 46.5730 0.2000 46.7730 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.096848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096848 LAYER M3 ;
    ANTENNAMAXAREACAR 32.48062 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.62056 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 40.76022 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.4930 0.0000 44.6930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.4930 0.0000 44.6930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.4930 0.0000 44.6930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.4930 0.0000 44.6930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.4930 0.0000 44.6930 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.298384 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.298384 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.7230 0.0000 42.9230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.7230 0.0000 42.9230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.7230 0.0000 42.9230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.7230 0.0000 42.9230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.7230 0.0000 42.9230 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 32.4540 87.6530 32.6540 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 32.4540 87.6530 32.6540 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 32.4540 87.6530 32.6540 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 32.4540 87.6530 32.6540 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 32.4540 87.6530 32.6540 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.135248 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.135248 LAYER M4 ;
    ANTENNAMAXAREACAR 59.04766 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 66.26283 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[3]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 48.6300 87.6530 48.8300 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 48.6300 87.6530 48.8300 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 48.6300 87.6530 48.8300 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 48.6300 87.6530 48.8300 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 48.6300 87.6530 48.8300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.2043 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.435826 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.435826 LAYER M2 ;
    ANTENNAMAXAREACAR 9.253289 LAYER M2 ;
    ANTENNAGATEAREA 0.6282 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 5.19262 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.19262 LAYER M3 ;
    ANTENNAMAXAREACAR 16.07485 LAYER M3 ;
    ANTENNAGATEAREA 0.6282 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 17.75931 LAYER M4 ;
    ANTENNAGATEAREA 0.6282 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.99947 LAYER M5 ;
    ANTENNAGATEAREA 0.6282 LAYER M6 ;
    ANTENNAGATEAREA 0.6282 LAYER M7 ;
    ANTENNAGATEAREA 0.6282 LAYER M8 ;
    ANTENNAGATEAREA 0.6282 LAYER M9 ;
    ANTENNAGATEAREA 0.6282 LAYER MRDL ;
  END SD

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 48.9700 87.6530 49.1700 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 48.9700 87.6530 49.1700 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 48.9700 87.6530 49.1700 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 48.9700 87.6530 49.1700 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 48.9700 87.6530 49.1700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.309528 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.309528 LAYER M2 ;
    ANTENNAMAXAREACAR 16.4589 LAYER M2 ;
    ANTENNAGATEAREA 0.0822 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 4.913532 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.913532 LAYER M3 ;
    ANTENNAMAXAREACAR 62.89865 LAYER M3 ;
    ANTENNAGATEAREA 0.0822 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 78.07346 LAYER M4 ;
    ANTENNAGATEAREA 0.0822 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 79.91259 LAYER M5 ;
    ANTENNAGATEAREA 0.0822 LAYER M6 ;
    ANTENNAGATEAREA 0.0822 LAYER M7 ;
    ANTENNAGATEAREA 0.0822 LAYER M8 ;
    ANTENNAGATEAREA 0.0822 LAYER M9 ;
    ANTENNAGATEAREA 0.0822 LAYER MRDL ;
  END DS1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 17.2900 87.6530 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 17.2900 87.6530 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 17.2900 87.6530 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 17.2900 87.6530 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 17.2900 87.6530 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30004 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30004 LAYER M4 ;
    ANTENNAMAXAREACAR 13.20148 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.63336 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 16.8310 87.6530 17.0310 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 16.8310 87.6530 17.0310 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 16.8310 87.6530 17.0310 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 16.8310 87.6530 17.0310 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 16.8310 87.6530 17.0310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.425149 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.425149 LAYER M4 ;
    ANTENNAMAXAREACAR 14.0694 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.21054 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 83.8260 58.8550 84.1250 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.7250 58.8550 85.0260 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9260 58.8550 2.2260 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.7250 58.8550 13.0250 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.0250 58.8550 1.3250 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8240 58.8550 12.1240 59.1550 ;
    END
    ANTENNADIFFAREA 11.07611 LAYER M5 ;
    ANTENNADIFFAREA 11.07611 LAYER M6 ;
    ANTENNADIFFAREA 11.07611 LAYER M7 ;
    ANTENNADIFFAREA 11.07611 LAYER M8 ;
    ANTENNADIFFAREA 11.07611 LAYER M9 ;
    ANTENNADIFFAREA 11.07611 LAYER MRDL ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 104.8005 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 104.8005 LAYER M5 ;
    ANTENNAMAXAREACAR 2644.257 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 5.9750 58.8550 6.2760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6750 58.8550 62.9760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8750 58.8550 7.1760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9750 58.8550 51.2740 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3750 58.8550 56.6750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4750 58.8550 55.7750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6750 58.8550 53.9750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5760 58.8550 54.8760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7750 58.8550 53.0750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8760 58.8550 52.1770 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0760 58.8550 50.3760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2750 58.8550 48.5750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4750 58.8550 46.7740 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6750 58.8550 44.9750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5760 58.8550 45.8760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1750 58.8550 49.4750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3760 58.8550 47.6770 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5760 58.8550 36.8750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0760 58.8550 41.3760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1750 58.8550 40.4750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9750 58.8550 42.2740 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7750 58.8550 44.0750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2750 58.8550 39.5750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4750 58.8550 37.7760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3750 58.8550 38.6760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8760 58.8550 43.1770 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1750 58.8550 85.4750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3750 58.8550 29.6750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0760 58.8550 86.3760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2760 58.8550 30.5760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1760 58.8550 31.4750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0760 58.8550 32.3750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7760 58.8550 35.0760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6760 58.8550 35.9750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8750 58.8550 34.1760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9750 58.8550 33.2760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8750 58.8550 79.1750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0750 58.8550 23.3750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9760 58.8550 78.2760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1760 58.8550 22.4760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6760 58.8550 80.9760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8760 58.8550 25.1760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5760 58.8550 81.8750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7760 58.8550 26.0750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3750 58.8550 83.6750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5750 58.8550 27.8750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2760 58.8550 84.5760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4760 58.8550 28.7760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4750 58.8550 82.7760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6750 58.8550 26.9760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7750 58.8550 80.0760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9750 58.8550 24.2760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.0760 58.8550 77.3760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2760 58.8550 21.5760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6750 58.8550 71.9750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8750 58.8550 16.1750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7760 58.8550 71.0760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9760 58.8550 15.2760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5760 58.8550 72.8750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7760 58.8550 17.0750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4750 58.8550 73.7750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6750 58.8550 17.9750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3750 58.8550 74.6760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5750 58.8550 18.8760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2750 58.8550 75.5760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4750 58.8550 19.7760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1750 58.8550 76.4760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3750 58.8550 20.6760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0760 58.8550 68.3760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2760 58.8550 12.5760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3760 58.8550 65.6750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5760 58.8550 9.8750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5760 58.8550 63.8760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7760 58.8550 8.0760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9760 58.8550 69.2750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1760 58.8550 13.4750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4760 58.8550 64.7750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6760 58.8550 8.9750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8750 58.8550 70.1750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0750 58.8550 14.3750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2750 58.8550 66.5760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4750 58.8550 10.7760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1750 58.8550 67.4760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3750 58.8550 11.6760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2760 58.8550 57.5750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4760 58.8550 1.7750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0750 58.8550 59.3750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2750 58.8550 3.5750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7750 58.8550 62.0760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3750 58.8550 2.6760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1750 58.8550 58.4760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0750 58.8550 5.3750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8750 58.8550 61.1750 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.1760 58.8550 4.4760 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9760 58.8550 60.2760 59.1550 ;
    END
  END VSS

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9900 0.0000 27.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9900 0.0000 27.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9900 0.0000 27.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9900 0.0000 27.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9900 0.0000 27.1900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6220 0.0000 25.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6220 0.0000 25.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6220 0.0000 25.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6220 0.0000 25.8220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2540 0.0010 24.4540 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2540 0.0010 24.4540 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2540 0.0000 24.4540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2540 0.0000 24.4540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2540 0.0000 24.4540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1514 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1514 LAYER M4 ;
    ANTENNAMAXAREACAR 69.58414 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1514 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1514 LAYER M5 ;
    ANTENNAMAXAREACAR 76.78907 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[15]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8860 0.0000 23.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8860 0.0000 23.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8860 0.0000 23.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8860 0.0000 23.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8860 0.0000 23.0860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.40786 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40786 LAYER M4 ;
    ANTENNAMAXAREACAR 13.59256 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.73374 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0894 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.31018 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.31018 LAYER M4 ;
    ANTENNAMAXAREACAR 6.388704 LAYER M4 ;
    ANTENNAGATEAREA 0.0894 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.084032 LAYER M5 ;
    ANTENNAGATEAREA 0.0894 LAYER M6 ;
    ANTENNAGATEAREA 0.0894 LAYER M7 ;
    ANTENNAGATEAREA 0.0894 LAYER M8 ;
    ANTENNAGATEAREA 0.0894 LAYER M9 ;
    ANTENNAGATEAREA 0.0894 LAYER MRDL ;
  END CE2

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 4.6250 58.8550 4.9260 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.5250 58.8550 5.8250 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.4250 58.8550 15.7260 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.3250 58.8550 16.6250 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.3250 58.8550 79.6250 59.1550 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.4260 58.8550 78.7260 59.1550 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 104.8014 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 104.8014 LAYER M5 ;
  END VDDL

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 52.6365 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 287.0016 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 287.0016 LAYER M2 ;
    ANTENNAMAXAREACAR 25.07252 LAYER M2 ;
    ANTENNAGATEAREA 55.8177 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 42.34068 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.34068 LAYER M3 ;
    ANTENNAMAXAREACAR 16.22651 LAYER M3 ;
    ANTENNAGATEAREA 55.8177 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 360.011 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 360.011 LAYER M4 ;
    ANTENNAMAXAREACAR 32.28083 LAYER M4 ;
    ANTENNAGATEAREA 55.8645 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 2867.268 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 2867.268 LAYER M5 ;
    ANTENNAMAXAREACAR 138.2991 LAYER M5 ;
    ANTENNAGATEAREA 55.8645 LAYER M6 ;
    ANTENNAGATEAREA 55.8645 LAYER M7 ;
    ANTENNAGATEAREA 55.8645 LAYER M8 ;
    ANTENNAGATEAREA 55.8645 LAYER M9 ;
    ANTENNAGATEAREA 55.8645 LAYER MRDL ;
  END WEB2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 52.1840 87.6530 52.3840 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 52.1840 87.6530 52.3840 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 52.1840 87.6530 52.3840 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 52.1840 87.6530 52.3840 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 52.1840 87.6530 52.3840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.298065 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.298065 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 30.09684 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 33.13903 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.18103 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 52.1720 0.2000 52.3720 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 52.1720 0.2000 52.3720 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 52.1720 0.2000 52.3720 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 52.1720 0.2000 52.3720 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 52.1720 0.2000 52.3720 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.234945 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.234945 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 28.37238 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.41469 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.45679 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 48.9580 0.2000 49.1580 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 48.9580 0.2000 49.1580 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 48.9580 0.2000 49.1580 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 48.9580 0.2000 49.1580 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 48.9580 0.2000 49.1580 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.246408 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.246408 LAYER M2 ;
    ANTENNAMAXAREACAR 13.49551 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.2326 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2326 LAYER M3 ;
    ANTENNAMAXAREACAR 29.71643 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 43.84799 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 47.16966 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5970 0.0000 20.7970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5970 0.0000 20.7970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5970 0.0000 20.7970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5970 0.0000 20.7970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5970 0.0000 20.7970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.2682 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.55632 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.55632 LAYER M2 ;
    ANTENNAMAXAREACAR 6.768853 LAYER M2 ;
    ANTENNAGATEAREA 0.2682 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 7.333657 LAYER M3 ;
    ANTENNAGATEAREA 0.2682 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.898423 LAYER M4 ;
    ANTENNAGATEAREA 0.2682 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.463151 LAYER M5 ;
    ANTENNAGATEAREA 0.2682 LAYER M6 ;
    ANTENNAGATEAREA 0.2682 LAYER M7 ;
    ANTENNAGATEAREA 0.2682 LAYER M8 ;
    ANTENNAGATEAREA 0.2682 LAYER M9 ;
    ANTENNAGATEAREA 0.2682 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8610 0.0000 67.0610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8610 0.0000 67.0610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8610 0.0000 67.0610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8610 0.0000 67.0610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8610 0.0000 67.0610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.2682 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56214 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56214 LAYER M2 ;
    ANTENNAMAXAREACAR 6.790553 LAYER M2 ;
    ANTENNAGATEAREA 0.2682 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 7.355355 LAYER M3 ;
    ANTENNAGATEAREA 0.2682 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.92012 LAYER M4 ;
    ANTENNAGATEAREA 0.2682 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.484847 LAYER M5 ;
    ANTENNAGATEAREA 0.2682 LAYER M6 ;
    ANTENNAGATEAREA 0.2682 LAYER M7 ;
    ANTENNAGATEAREA 0.2682 LAYER M8 ;
    ANTENNAGATEAREA 0.2682 LAYER M9 ;
    ANTENNAGATEAREA 0.2682 LAYER MRDL ;
  END OEB1

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.3840 0.0000 53.5840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.3840 0.0000 53.5840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.3840 0.0000 53.5840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.3840 0.0000 53.5840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.3840 0.0000 53.5840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.0160 0.0000 52.2160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.0160 0.0000 52.2160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.0160 0.0000 52.2160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.0160 0.0000 52.2160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.0160 0.0000 52.2160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.6480 0.0000 50.8480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.6480 0.0000 50.8480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.6480 0.0000 50.8480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.6480 0.0000 50.8480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.6480 0.0000 50.8480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.2800 0.0000 49.4800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.2800 0.0000 49.4800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.2800 0.0000 49.4800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.2800 0.0000 49.4800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.2800 0.0000 49.4800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.9120 0.0000 48.1120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.9120 0.0000 48.1120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.9120 0.0000 48.1120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.9120 0.0000 48.1120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.9120 0.0000 48.1120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.5440 0.0000 46.7440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.5440 0.0000 46.7440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.5440 0.0000 46.7440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.5440 0.0000 46.7440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.5440 0.0000 46.7440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.1760 0.0000 45.3760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.1760 0.0000 45.3760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.1760 0.0000 45.3760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.1760 0.0000 45.3760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.1760 0.0000 45.3760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.4060 0.0000 43.6060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.4060 0.0000 43.6060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.4060 0.0000 43.6060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.4060 0.0000 43.6060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.4060 0.0000 43.6060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0380 0.0000 42.2380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0380 0.0000 42.2380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0380 0.0000 42.2380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0380 0.0000 42.2380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0380 0.0000 42.2380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6700 0.0000 40.8700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6700 0.0000 40.8700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6700 0.0000 40.8700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6700 0.0000 40.8700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6700 0.0000 40.8700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.3020 0.0000 39.5020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.3020 0.0000 39.5020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.3020 0.0000 39.5020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.3020 0.0000 39.5020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.3020 0.0000 39.5020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9340 0.0000 38.1340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9340 0.0000 38.1340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9340 0.0000 38.1340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9340 0.0000 38.1340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9340 0.0000 38.1340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5660 0.0000 36.7660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5660 0.0000 36.7660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5660 0.0000 36.7660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5660 0.0000 36.7660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5660 0.0000 36.7660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1980 0.0000 35.3980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1980 0.0000 35.3980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1980 0.0000 35.3980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1980 0.0000 35.3980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1980 0.0000 35.3980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8300 0.0000 34.0300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8300 0.0000 34.0300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8300 0.0000 34.0300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8300 0.0000 34.0300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8300 0.0000 34.0300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4620 0.0000 32.6620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4620 0.0000 32.6620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4620 0.0000 32.6620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4620 0.0000 32.6620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4620 0.0000 32.6620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0940 0.0000 31.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0940 0.0000 31.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0940 0.0000 31.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0940 0.0000 31.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0940 0.0000 31.2940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7260 0.0000 29.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7260 0.0000 29.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7260 0.0000 29.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7260 0.0000 29.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7260 0.0000 29.9260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3580 0.0000 28.5580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3580 0.0000 28.5580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3580 0.0000 28.5580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3580 0.0000 28.5580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3580 0.0000 28.5580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.7010 0.0000 52.9010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.7010 0.0000 52.9010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.7010 0.0000 52.9010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.7010 0.0000 52.9010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.7010 0.0000 52.9010 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4370 0.0000 55.6370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4370 0.0000 55.6370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4370 0.0000 55.6370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4370 0.0000 55.6370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4370 0.0000 55.6370 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.0690 0.0000 54.2690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.0690 0.0000 54.2690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.0690 0.0000 54.2690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.0690 0.0000 54.2690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.0690 0.0000 54.2690 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.1730 0.0000 58.3730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.1730 0.0000 58.3730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.1730 0.0000 58.3730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.1730 0.0000 58.3730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.1730 0.0000 58.3730 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.5410 0.0000 59.7410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.5410 0.0000 59.7410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.5410 0.0000 59.7410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.5410 0.0000 59.7410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.5410 0.0000 59.7410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[0]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.9090 0.0000 61.1090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.9090 0.0000 61.1090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.9090 0.0000 61.1090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.9090 0.0000 61.1090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.9090 0.0000 61.1090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[14]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.2770 0.0000 62.4770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.2770 0.0000 62.4770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.2770 0.0000 62.4770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.2770 0.0000 62.4770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.2770 0.0000 62.4770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.6450 0.0000 63.8450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.6450 0.0000 63.8450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.6450 0.0000 63.8450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.6450 0.0000 63.8450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.6450 0.0000 63.8450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[8]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.0130 0.0000 65.2130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.0130 0.0000 65.2130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.0130 0.0000 65.2130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.0130 0.0000 65.2130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.0130 0.0000 65.2130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[10]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.3810 0.0000 66.5810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.3810 0.0000 66.5810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.3810 0.0000 66.5810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.3810 0.0000 66.5810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.3810 0.0000 66.5810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[3]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.6960 0.0000 65.8960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.6960 0.0000 65.8960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.6960 0.0000 65.8960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.6960 0.0000 65.8960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6960 0.0000 65.8960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.3280 0.0000 64.5280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.3280 0.0000 64.5280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.3280 0.0000 64.5280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.3280 0.0000 64.5280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.3280 0.0000 64.5280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.9600 0.0000 63.1600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.9600 0.0000 63.1600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.9600 0.0000 63.1600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.9600 0.0000 63.1600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.9600 0.0000 63.1600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.5920 0.0000 61.7920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.5920 0.0000 61.7920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.5920 0.0000 61.7920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.5920 0.0000 61.7920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.5920 0.0000 61.7920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.2240 0.0000 60.4240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.2240 0.0000 60.4240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.2240 0.0000 60.4240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.2240 0.0000 60.4240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.2240 0.0000 60.4240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.8560 0.0000 59.0560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.8560 0.0000 59.0560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.8560 0.0000 59.0560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.8560 0.0000 59.0560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.8560 0.0000 59.0560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.4880 0.0000 57.6880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.4880 0.0000 57.6880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.4880 0.0000 57.6880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.4880 0.0000 57.6880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.4880 0.0000 57.6880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7520 0.0000 54.9520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7520 0.0000 54.9520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7520 0.0000 54.9520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7520 0.0000 54.9520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7520 0.0000 54.9520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.3550 0.0000 41.5550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.3550 0.0000 41.5550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.3550 0.0000 41.5550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.3550 0.0000 41.5550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.3550 0.0000 41.5550 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9870 0.0000 40.1870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9870 0.0000 40.1870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9870 0.0000 40.1870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9870 0.0000 40.1870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9870 0.0000 40.1870 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.6190 0.0000 38.8190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.6190 0.0000 38.8190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.6190 0.0000 38.8190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.6190 0.0000 38.8190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.6190 0.0000 38.8190 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.2510 0.0000 37.4510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.2510 0.0000 37.4510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.2510 0.0000 37.4510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.2510 0.0000 37.4510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.2510 0.0000 37.4510 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8830 0.0000 36.0830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8830 0.0000 36.0830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8830 0.0000 36.0830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8830 0.0000 36.0830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8830 0.0000 36.0830 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.5150 0.0000 34.7150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.5150 0.0000 34.7150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.5150 0.0000 34.7150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.5150 0.0000 34.7150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.5150 0.0000 34.7150 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1470 0.0000 33.3470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1470 0.0000 33.3470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1470 0.0000 33.3470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1470 0.0000 33.3470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1470 0.0000 33.3470 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7790 0.0000 31.9790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7790 0.0000 31.9790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7790 0.0000 31.9790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7790 0.0000 31.9790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7790 0.0000 31.9790 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.4110 0.0000 30.6110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.4110 0.0000 30.6110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.4110 0.0000 30.6110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.4110 0.0000 30.6110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.4110 0.0000 30.6110 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.0430 0.0000 29.2430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.0430 0.0000 29.2430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.0430 0.0000 29.2430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.0430 0.0000 29.2430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.0430 0.0000 29.2430 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[11]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6750 0.0000 27.8750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6750 0.0000 27.8750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6750 0.0000 27.8750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6750 0.0000 27.8750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6750 0.0000 27.8750 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[4]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.3070 0.0000 26.5070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.3070 0.0000 26.5070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.3070 0.0000 26.5070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.3070 0.0000 26.5070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.3070 0.0000 26.5070 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[2]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.1200 0.0000 56.3200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.1200 0.0000 56.3200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.1200 0.0000 56.3200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.1200 0.0000 56.3200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.1200 0.0000 56.3200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.8050 0.0000 57.0050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.8050 0.0000 57.0050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.8050 0.0000 57.0050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.8050 0.0000 57.0050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.8050 0.0000 57.0050 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.8610 0.0000 46.0610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.8610 0.0000 46.0610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.8610 0.0000 46.0610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.8610 0.0000 46.0610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.8610 0.0000 46.0610 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.2290 0.0000 47.4290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.2290 0.0000 47.4290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.2290 0.0000 47.4290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.2290 0.0000 47.4290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.2290 0.0000 47.4290 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.5970 0.0000 48.7970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.5970 0.0000 48.7970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.5970 0.0000 48.7970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.5970 0.0000 48.7970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.5970 0.0000 48.7970 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.9650 0.0000 50.1650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.9650 0.0000 50.1650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.9650 0.0000 50.1650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.9650 0.0000 50.1650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.9650 0.0000 50.1650 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.3330 0.0000 51.5330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.3330 0.0000 51.5330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.3330 0.0000 51.5330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.3330 0.0000 51.5330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.3330 0.0000 51.5330 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 46.5840 87.6530 46.7840 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 46.5840 87.6530 46.7840 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 46.5840 87.6530 46.7840 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 46.5840 87.6530 46.7840 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 46.5840 87.6530 46.7840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.096188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096188 LAYER M3 ;
    ANTENNAMAXAREACAR 32.46259 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.60252 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 40.74219 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 39.2840 87.6530 39.4840 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 39.2840 87.6530 39.4840 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 39.2840 87.6530 39.4840 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 39.2840 87.6530 39.4840 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 39.2840 87.6530 39.4840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.096188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096188 LAYER M3 ;
    ANTENNAMAXAREACAR 32.46259 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.60252 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 40.74219 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 37.7610 87.6530 37.9610 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 37.7610 87.6530 37.9610 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 37.7610 87.6530 37.9610 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 37.7610 87.6530 37.9610 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 37.7610 87.6530 37.9610 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.096188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096188 LAYER M3 ;
    ANTENNAMAXAREACAR 32.46259 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.60252 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 40.74219 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[2]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4530 9.8210 87.6530 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4530 9.8210 87.6530 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4530 9.8210 87.6530 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4530 9.8210 87.6530 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4530 9.8210 87.6530 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
  END WEB1

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.9390 0.0000 25.1390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.9390 0.0000 25.1390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.9390 0.0000 25.1390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.9390 0.0000 25.1390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.9390 0.0000 25.1390 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[15]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5710 0.0000 23.7710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5710 0.0000 23.7710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5710 0.0000 23.7710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5710 0.0000 23.7710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5710 0.0000 23.7710 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[6]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.4890 0.2000 32.6890 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 32.4890 0.2000 32.6890 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 32.4890 0.2000 32.6890 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.4890 0.2000 32.6890 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 32.4890 0.2000 32.6890 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.134288 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.134288 LAYER M4 ;
    ANTENNAMAXAREACAR 59.1957 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 66.41084 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 37.7580 0.2000 37.9580 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 37.7580 0.2000 37.9580 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 37.7580 0.2000 37.9580 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 37.7580 0.2000 37.9580 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 37.7580 0.2000 37.9580 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.096848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096848 LAYER M3 ;
    ANTENNAMAXAREACAR 32.48062 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.62056 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 40.76022 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 39.2760 0.2000 39.4760 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 39.2760 0.2000 39.4760 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 39.2760 0.2000 39.4760 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 39.2760 0.2000 39.4760 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 39.2760 0.2000 39.4760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.096848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096848 LAYER M3 ;
    ANTENNAMAXAREACAR 32.48062 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 36.62056 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 40.76022 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]
  OBS
    LAYER M1 ;
      RECT 86.8530 38.5610 87.6530 38.5750 ;
      RECT 0.8000 38.6840 86.8530 40.0760 ;
      RECT 0.8000 38.6760 87.6530 38.6840 ;
      RECT 0.0000 38.5580 0.8000 38.5750 ;
      RECT 0.0000 47.3730 0.8000 48.3580 ;
      RECT 0.0000 0.0000 19.9970 0.8000 ;
      RECT 0.8000 31.8890 86.8530 33.2540 ;
      RECT 0.8000 38.5610 86.8530 38.6760 ;
      RECT 0.8000 38.5580 86.8530 38.5610 ;
      RECT 0.0000 31.8540 86.8530 31.8890 ;
      RECT 0.0000 0.0000 19.9970 9.2210 ;
      RECT 0.0000 18.1680 86.8530 31.8890 ;
      RECT 0.0000 18.1680 86.8530 31.8890 ;
      RECT 0.0000 18.1680 86.8530 31.8890 ;
      RECT 0.0000 18.1680 87.6530 31.8540 ;
      RECT 0.8000 18.1680 86.8530 33.2540 ;
      RECT 0.8000 18.1680 86.8530 33.2540 ;
      RECT 0.8000 18.1680 86.8530 33.2540 ;
      RECT 0.0000 16.2310 86.8530 16.2340 ;
      RECT 0.0000 10.6210 86.8530 16.2340 ;
      RECT 0.0000 10.6210 86.8530 16.2340 ;
      RECT 0.0000 10.6210 86.8530 16.2340 ;
      RECT 0.0000 10.6210 87.6530 16.2310 ;
      RECT 0.8000 18.0900 87.6530 31.8540 ;
      RECT 0.8000 18.0900 87.6530 31.8540 ;
      RECT 0.8000 18.0900 87.6530 31.8540 ;
      RECT 0.8000 18.0900 87.6530 18.1680 ;
      RECT 0.8000 16.2340 86.8530 18.0900 ;
      RECT 0.8000 10.6210 86.8530 18.0900 ;
      RECT 0.8000 10.6210 86.8530 18.0900 ;
      RECT 0.8000 10.6210 86.8530 18.0900 ;
      RECT 0.8000 9.2210 86.8530 16.2310 ;
      RECT 0.8000 9.2210 86.8530 10.6210 ;
      RECT 0.0000 0.8000 87.6530 9.2210 ;
      RECT 67.6610 0.0000 87.6530 9.2210 ;
      RECT 67.6610 0.0000 87.6530 0.8000 ;
      RECT 0.0000 52.9840 87.6530 59.1550 ;
      RECT 0.8000 48.0300 86.8530 48.3580 ;
      RECT 0.8000 49.7700 86.8530 59.1550 ;
      RECT 0.8000 49.7700 86.8530 59.1550 ;
      RECT 0.8000 49.7700 86.8530 59.1550 ;
      RECT 0.8000 48.3580 86.8530 59.1550 ;
      RECT 0.8000 48.3580 86.8530 59.1550 ;
      RECT 0.8000 48.3580 86.8530 59.1550 ;
      RECT 0.0000 40.0840 87.6530 45.9730 ;
      RECT 0.8000 45.9840 86.8530 52.9840 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 52.9720 ;
      RECT 0.8000 45.9840 86.8530 51.5840 ;
      RECT 0.8000 45.9840 86.8530 51.5840 ;
      RECT 0.8000 45.9840 86.8530 49.7700 ;
      RECT 0.8000 45.9840 86.8530 49.7700 ;
      RECT 0.8000 40.0840 86.8530 49.7700 ;
      RECT 0.8000 40.0840 86.8530 49.7700 ;
      RECT 0.8000 40.0840 86.8530 49.7700 ;
      RECT 0.8000 40.0840 86.8530 49.7700 ;
      RECT 0.8000 40.0840 86.8530 49.7580 ;
      RECT 0.8000 40.0840 86.8530 49.7580 ;
      RECT 0.8000 40.0840 86.8530 49.7580 ;
      RECT 0.8000 40.0840 86.8530 49.7580 ;
      RECT 0.8000 40.0840 86.8530 49.7580 ;
      RECT 0.8000 40.0840 86.8530 49.7580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.8000 40.0840 86.8530 48.3580 ;
      RECT 0.0000 33.2890 87.6530 37.1580 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2890 86.8530 38.6840 ;
      RECT 0.8000 33.2540 87.6530 37.1580 ;
      RECT 0.8000 33.2540 87.6530 37.1580 ;
      RECT 0.8000 33.2540 87.6530 37.1580 ;
      RECT 0.8000 33.2540 87.6530 33.2890 ;
      RECT 86.8530 47.3840 87.6530 48.0300 ;
      RECT 21.3970 0.0000 22.2860 0.8000 ;
      RECT 0.0000 49.7580 1.5010 51.5720 ;
      RECT 0.0000 40.0760 86.8530 43.0770 ;
      RECT 0.0000 52.9720 3.0010 52.9840 ;
      RECT 86.1520 49.7700 87.6530 51.5840 ;
      RECT 84.6520 45.9730 87.6530 45.9840 ;
      RECT 84.6520 37.1580 87.6530 37.1610 ;
      RECT 0.0000 38.5750 87.6530 38.6760 ;
    LAYER PO ;
      RECT 0.0000 0.0000 87.6530 59.1550 ;
    LAYER M3 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 87.6530 31.7540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.0000 16.1310 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 87.6530 16.1310 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 18.2680 ;
      RECT 0.9000 16.1340 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 9.1210 86.7530 10.7210 ;
      RECT 0.9000 0.9000 86.7530 10.7210 ;
      RECT 21.4970 0.0000 22.1860 0.9000 ;
      RECT 0.0000 47.4730 0.9000 48.2580 ;
      RECT 0.0000 49.8580 1.5010 51.4720 ;
      RECT 86.1520 49.8700 87.6530 51.4840 ;
      RECT 86.7530 47.4840 87.6530 47.9300 ;
      RECT 0.0000 40.1760 86.7530 40.1840 ;
      RECT 0.9000 37.0610 86.7530 40.1760 ;
      RECT 0.0000 0.0000 19.8970 9.1210 ;
      RECT 0.0000 0.9000 87.6530 9.1210 ;
      RECT 0.0000 0.0000 19.8970 0.9000 ;
      RECT 67.7610 0.0000 87.6530 9.1210 ;
      RECT 67.7610 0.0000 87.6530 0.9000 ;
      RECT 0.0000 53.0840 87.6530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 53.0840 ;
      RECT 0.9000 51.4840 86.7530 53.0720 ;
      RECT 0.0000 40.1840 87.6530 45.8730 ;
      RECT 0.0000 40.1760 86.7530 45.8730 ;
      RECT 0.9000 49.8700 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 53.0840 ;
      RECT 0.9000 45.8840 86.7530 53.0720 ;
      RECT 0.9000 45.8840 86.7530 53.0720 ;
      RECT 0.9000 45.8730 86.7530 53.0720 ;
      RECT 0.9000 51.4720 86.7530 51.4840 ;
      RECT 0.9000 48.2580 86.7530 51.4840 ;
      RECT 0.9000 48.2580 86.7530 51.4840 ;
      RECT 0.9000 45.8840 86.7530 51.4840 ;
      RECT 0.9000 45.8840 86.7530 51.4840 ;
      RECT 0.9000 45.8730 86.7530 51.4840 ;
      RECT 0.9000 49.8700 86.7530 51.4720 ;
      RECT 0.9000 48.2580 86.7530 51.4720 ;
      RECT 0.9000 48.2580 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 49.8580 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 48.2580 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 47.9300 86.7530 48.2580 ;
      RECT 0.9000 47.4840 86.7530 47.9300 ;
      RECT 0.9000 47.4730 86.7530 47.4840 ;
      RECT 0.9000 45.8840 86.7530 47.4730 ;
      RECT 0.9000 45.8730 87.6530 45.8840 ;
      RECT 0.9000 37.0610 86.7530 45.8730 ;
      RECT 0.0000 33.3890 87.6530 37.0580 ;
      RECT 0.9000 33.3890 86.7530 40.1760 ;
      RECT 0.9000 37.0580 87.6530 37.0610 ;
      RECT 0.9000 33.3890 87.6530 37.0610 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 33.3890 ;
      RECT 0.9000 31.7890 86.7530 33.3540 ;
      RECT 0.0000 31.7540 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
    LAYER M2 ;
      RECT 86.7530 47.4840 87.6530 47.9300 ;
      RECT 21.4970 0.0000 22.1860 0.9000 ;
      RECT 0.0000 49.8580 1.5010 51.4720 ;
      RECT 86.1520 49.8700 87.6530 51.4840 ;
      RECT 0.0000 47.4730 0.9000 48.2580 ;
      RECT 0.0000 40.1760 86.7530 40.1840 ;
      RECT 0.9000 37.0610 86.7530 40.1760 ;
      RECT 0.0000 0.0000 19.8970 9.1210 ;
      RECT 0.0000 0.9000 87.6530 9.1210 ;
      RECT 0.0000 0.0000 19.8970 0.9000 ;
      RECT 67.7610 0.0000 87.6530 9.1210 ;
      RECT 67.7610 0.0000 87.6530 0.9000 ;
      RECT 0.0000 53.0840 87.6530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 59.1550 ;
      RECT 0.0000 53.0720 86.7530 53.0840 ;
      RECT 0.9000 51.4840 86.7530 53.0720 ;
      RECT 0.0000 40.1840 87.6530 45.8730 ;
      RECT 0.0000 40.1760 86.7530 45.8730 ;
      RECT 0.9000 49.8700 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 53.0840 ;
      RECT 0.9000 45.8840 86.7530 53.0720 ;
      RECT 0.9000 45.8840 86.7530 53.0720 ;
      RECT 0.9000 45.8730 86.7530 53.0720 ;
      RECT 0.9000 51.4720 86.7530 51.4840 ;
      RECT 0.9000 48.2580 86.7530 51.4840 ;
      RECT 0.9000 48.2580 86.7530 51.4840 ;
      RECT 0.9000 45.8840 86.7530 51.4840 ;
      RECT 0.9000 45.8840 86.7530 51.4840 ;
      RECT 0.9000 45.8730 86.7530 51.4840 ;
      RECT 0.9000 49.8700 86.7530 51.4720 ;
      RECT 0.9000 48.2580 86.7530 51.4720 ;
      RECT 0.9000 48.2580 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 45.8730 86.7530 51.4720 ;
      RECT 0.9000 49.8580 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8840 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 45.8730 86.7530 49.8700 ;
      RECT 0.9000 48.2580 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 47.9300 86.7530 48.2580 ;
      RECT 0.9000 47.4840 86.7530 47.9300 ;
      RECT 0.9000 47.4730 86.7530 47.4840 ;
      RECT 0.9000 45.8840 86.7530 47.4730 ;
      RECT 0.9000 45.8730 87.6530 45.8840 ;
      RECT 0.9000 37.0610 86.7530 45.8730 ;
      RECT 0.0000 33.3890 87.6530 37.0580 ;
      RECT 0.9000 33.3890 86.7530 40.1760 ;
      RECT 0.9000 37.0580 87.6530 37.0610 ;
      RECT 0.9000 33.3890 87.6530 37.0610 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 33.3890 ;
      RECT 0.9000 31.7890 86.7530 33.3540 ;
      RECT 0.0000 31.7540 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 87.6530 31.7540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.0000 16.1310 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 87.6530 16.1310 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 18.2680 ;
      RECT 0.9000 16.1340 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 9.1210 86.7530 10.7210 ;
      RECT 0.9000 0.9000 86.7530 10.7210 ;
    LAYER M4 ;
      RECT 0.0000 31.7540 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 87.6530 31.7540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 18.2680 ;
      RECT 0.9000 16.1340 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.0000 0.9010 87.6530 9.1210 ;
      RECT 0.9000 9.1210 86.7530 16.1310 ;
      RECT 0.9000 9.1210 86.7530 10.7210 ;
      RECT 25.1540 0.9000 87.6530 9.1210 ;
      RECT 25.1540 0.9000 87.6530 9.1210 ;
      RECT 25.1540 0.9000 87.6530 9.1210 ;
      RECT 25.1540 0.9000 87.6530 0.9010 ;
      RECT 67.7610 0.0000 87.6530 9.1210 ;
      RECT 67.7610 0.0000 87.6530 9.1210 ;
      RECT 67.7610 0.0000 87.6530 0.9000 ;
      RECT 0.9000 47.9300 86.7530 48.2580 ;
      RECT 0.9000 47.4840 86.7530 47.9300 ;
      RECT 0.0000 53.0840 87.6530 59.1550 ;
      RECT 0.9000 49.8700 86.7530 59.1550 ;
      RECT 0.9000 49.8700 86.7530 59.1550 ;
      RECT 0.9000 49.8700 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 59.1550 ;
      RECT 0.9000 48.2580 86.7530 59.1550 ;
      RECT 0.9000 47.9300 86.7530 53.0840 ;
      RECT 0.9000 47.9300 86.7530 53.0720 ;
      RECT 0.9000 47.9300 86.7530 53.0720 ;
      RECT 0.9000 47.9300 86.7530 53.0720 ;
      RECT 0.9000 47.9300 86.7530 53.0720 ;
      RECT 0.9000 47.9300 86.7530 53.0720 ;
      RECT 0.9000 47.9300 86.7530 51.4720 ;
      RECT 0.9000 47.9300 86.7530 51.4720 ;
      RECT 0.9000 47.9300 86.7530 51.4720 ;
      RECT 0.9000 47.9300 86.7530 51.4720 ;
      RECT 0.0000 40.1840 87.6530 45.8730 ;
      RECT 0.0000 40.1760 86.7530 45.8730 ;
      RECT 0.0000 40.1760 86.7530 40.1840 ;
      RECT 0.9000 37.0610 86.7530 45.8730 ;
      RECT 21.4970 0.0000 22.1860 0.9000 ;
      RECT 0.0000 47.9300 86.7530 48.2580 ;
      RECT 0.0000 47.4840 87.6530 47.9300 ;
      RECT 0.0000 47.4730 86.7530 47.4840 ;
      RECT 0.0000 49.8580 1.5010 51.4720 ;
      RECT 0.0000 53.0720 3.0010 53.0840 ;
      RECT 0.9000 42.8830 87.6530 45.8840 ;
      RECT 0.9000 48.2580 86.7530 48.9740 ;
      RECT 0.9000 45.8840 86.7530 47.4730 ;
      RECT 86.1520 49.8700 87.6530 51.4840 ;
      RECT 0.0000 0.0000 19.8970 0.9000 ;
      RECT 0.0000 0.9000 23.5540 0.9010 ;
      RECT 0.0000 0.0000 19.8970 9.1210 ;
      RECT 0.0000 0.0000 19.8970 9.1210 ;
      RECT 0.0000 0.9000 23.5540 9.1210 ;
      RECT 0.0000 0.9000 23.5540 9.1210 ;
      RECT 0.0000 0.9000 23.5540 9.1210 ;
      RECT 0.9000 37.0610 86.7530 40.1760 ;
      RECT 0.0000 33.3890 87.6530 37.0580 ;
      RECT 0.9000 33.3890 86.7530 40.1760 ;
      RECT 0.9000 37.0580 87.6530 37.0610 ;
      RECT 0.9000 33.3890 87.6530 37.0610 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 33.3890 ;
      RECT 0.9000 31.7890 86.7530 33.3540 ;
      RECT 0.0000 16.1310 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 87.6530 16.1310 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 87.6530 59.1550 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 87.6530 59.1550 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 87.6530 59.1550 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 87.6530 59.1550 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 87.6530 59.1550 ;
    LAYER M5 ;
      RECT 0.0000 58.1550 0.3250 59.1550 ;
      RECT 21.4970 0.0000 22.1860 0.9000 ;
      RECT 87.0760 58.1550 87.6530 59.1550 ;
      RECT 0.0000 47.4730 0.9000 48.2580 ;
      RECT 0.0000 53.0720 3.0010 53.0840 ;
      RECT 0.0000 49.8580 1.5010 51.4720 ;
      RECT 0.9000 42.8830 87.6530 45.8840 ;
      RECT 86.1520 49.8700 87.6530 51.4840 ;
      RECT 86.7530 47.4840 87.6530 47.9300 ;
      RECT 0.0000 0.0000 19.8970 0.9000 ;
      RECT 0.0000 0.9000 23.5540 0.9010 ;
      RECT 0.0000 0.0000 19.8970 9.1210 ;
      RECT 0.0000 0.0000 19.8970 9.1210 ;
      RECT 0.0000 0.9000 23.5540 9.1210 ;
      RECT 0.0000 0.9000 23.5540 9.1210 ;
      RECT 0.0000 0.9000 23.5540 9.1210 ;
      RECT 0.9000 31.7890 86.7530 33.3540 ;
      RECT 0.0000 31.7540 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 86.7530 31.7890 ;
      RECT 0.0000 18.2680 87.6530 31.7540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.9000 18.2680 86.7530 33.3540 ;
      RECT 0.0000 33.3890 87.6530 37.0580 ;
      RECT 0.9000 37.0610 86.7530 40.1760 ;
      RECT 0.9000 33.3890 86.7530 40.1760 ;
      RECT 0.9000 37.0580 87.6530 37.0610 ;
      RECT 0.9000 33.3890 87.6530 37.0610 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 37.0580 ;
      RECT 0.9000 33.3540 87.6530 33.3890 ;
      RECT 0.0000 16.1310 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 86.7530 16.1340 ;
      RECT 0.0000 10.7210 87.6530 16.1310 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 31.7540 ;
      RECT 0.9000 18.1900 87.6530 18.2680 ;
      RECT 0.9000 16.1340 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.9000 10.7210 86.7530 18.1900 ;
      RECT 0.0000 0.9010 87.6530 9.1210 ;
      RECT 0.9000 9.1210 86.7530 16.1310 ;
      RECT 0.9000 9.1210 86.7530 10.7210 ;
      RECT 25.1540 0.9000 87.6530 9.1210 ;
      RECT 25.1540 0.9000 87.6530 9.1210 ;
      RECT 25.1540 0.9000 87.6530 9.1210 ;
      RECT 25.1540 0.9000 87.6530 0.9010 ;
      RECT 67.7610 0.0000 87.6530 9.1210 ;
      RECT 67.7610 0.0000 87.6530 9.1210 ;
      RECT 67.7610 0.0000 87.6530 0.9000 ;
      RECT 0.9000 47.9300 86.7530 48.2580 ;
      RECT 0.0000 53.0840 87.6530 58.1550 ;
      RECT 0.0000 40.1840 87.6530 45.8730 ;
      RECT 0.0000 40.1760 86.7530 45.8730 ;
      RECT 0.0000 40.1760 86.7530 40.1840 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 45.8840 86.7530 49.8580 ;
      RECT 0.9000 37.0610 86.7530 45.8730 ;
      RECT 0.9000 49.8700 86.7530 58.1550 ;
      RECT 0.9000 49.8700 86.7530 58.1550 ;
      RECT 0.9000 49.8700 86.7530 58.1550 ;
      RECT 0.9000 49.8700 86.7530 58.1550 ;
      RECT 0.9000 48.2580 86.7530 58.1550 ;
      RECT 0.9000 48.2580 86.7530 58.1550 ;
      RECT 0.9000 48.2580 86.7530 58.1550 ;
      RECT 0.9000 48.2580 86.7530 53.0840 ;
      RECT 0.9000 48.2580 86.7530 53.0840 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
      RECT 0.9000 45.8840 86.7530 51.4720 ;
  END
END SRAMLP2RW16x16

MACRO SRAMLP2RW16x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 131.406 BY 68.044 ;
  SYMMETRY X Y R90 ;

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[30]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.5440 0.0000 74.7440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.5440 0.0000 74.7440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.5440 0.0000 74.7440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.5440 0.0000 74.7440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.5440 0.0000 74.7440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.8080 0.0000 72.0080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.8080 0.0000 72.0080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.8080 0.0000 72.0080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.8080 0.0000 72.0080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.8080 0.0000 72.0080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[19]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.1760 0.0000 73.3760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.1760 0.0000 73.3760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.1760 0.0000 73.3760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.1760 0.0000 73.3760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.1760 0.0000 73.3760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[30]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.7050 0.0000 67.9050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.7040 0.0000 67.9040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.7040 0.0000 67.9040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.7040 0.0000 67.9040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.7040 0.0000 67.9040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.0720 0.0000 69.2720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.0720 0.0000 69.2720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.0720 0.0000 69.2720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.0720 0.0000 69.2720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.0720 0.0000 69.2720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.7290 0.0000 65.9290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.7290 0.0000 65.9290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.7290 0.0000 65.9290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.7290 0.0000 65.9290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.7290 0.0000 65.9290 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.265908 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.265908 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.4400 0.0000 70.6400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.4400 0.0000 70.6400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.4400 0.0000 70.6400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.4400 0.0000 70.6400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4400 0.0000 70.6400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[14]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[21]

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 126.1040 67.7440 126.4030 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.0040 67.7440 127.3030 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.5080 67.7440 14.8080 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.4090 67.7440 15.7090 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.7080 67.7440 4.0080 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.6090 67.7440 4.9080 68.0440 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 120.6642 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 120.6642 LAYER M5 ;
  END VDDL

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.3280 0.0000 92.5280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.3280 0.0000 92.5280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.3280 0.0000 92.5280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.3280 0.0000 92.5280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.3280 0.0000 92.5280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[21]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6960 0.0000 93.8960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6960 0.0000 93.8960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6960 0.0000 93.8960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6960 0.0000 93.8960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6960 0.0000 93.8960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.9600 0.0000 91.1600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.9600 0.0000 91.1600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.9600 0.0000 91.1600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.9600 0.0000 91.1600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.9600 0.0000 91.1600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[29]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.1200 0.0000 84.3200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.1200 0.0000 84.3200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.1200 0.0000 84.3200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.1200 0.0000 84.3200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.1200 0.0000 84.3200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[23]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.29355 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29355 LAYER M3 ;
    ANTENNAMAXAREACAR 62.84588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 70.06078 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.27521 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[26]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.4880 0.0000 85.6880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.4880 0.0000 85.6880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.4880 0.0000 85.6880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.4880 0.0000 85.6880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.4880 0.0000 85.6880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.8560 0.0000 87.0560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.8560 0.0000 87.0560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.8560 0.0000 87.0560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.8560 0.0000 87.0560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.8560 0.0000 87.0560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[31]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.8300 -0.0020 85.0300 0.1980 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.8300 -0.0020 85.0300 0.1980 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.8300 -0.0020 85.0300 0.1980 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.8300 -0.0020 85.0300 0.1980 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.8300 -0.0020 85.0300 0.1980 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28848 LAYER M3 ;
    ANTENNAMAXAREACAR 62.60445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81937 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.03381 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[31]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[22]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.2240 0.0000 88.4240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.2240 0.0000 88.4240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.2240 0.0000 88.4240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.2240 0.0000 88.4240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.2240 0.0000 88.4240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[26]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[28]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.9120 0.0000 76.1120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.9120 0.0000 76.1120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.9120 0.0000 76.1120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.9120 0.0000 76.1120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.9120 0.0000 76.1120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.2800 0.0000 77.4800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.2800 0.0000 77.4800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.2800 0.0000 77.4800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.2800 0.0000 77.4800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.2800 0.0000 77.4800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.0080 0.0000 106.2080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.0080 0.0000 106.2080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.0080 0.0000 106.2080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.0080 0.0000 106.2080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.0080 0.0000 106.2080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[18]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[17]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.9040 0.0000 102.1040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.9040 0.0000 102.1040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.9040 0.0000 102.1040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.9040 0.0000 102.1040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.9040 0.0000 102.1040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[17]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.6400 0.0000 104.8400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.6400 0.0000 104.8400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.6400 0.0000 104.8400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.6400 0.0000 104.8400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.6400 0.0000 104.8400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[9]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.1680 0.0000 99.3680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.1680 0.0000 99.3680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.1680 0.0000 99.3680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.1680 0.0000 99.3680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.1680 0.0000 99.3680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[20]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[24]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.4320 0.0000 96.6320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.4320 0.0000 96.6320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.4320 0.0000 96.6320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.4320 0.0000 96.6320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.4320 0.0000 96.6320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[20]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.8010 0.0000 98.0010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.8010 0.0000 98.0010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.8010 0.0000 98.0010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.8010 0.0000 98.0010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.8010 0.0000 98.0010 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[24]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[27]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.0640 0.0000 95.2640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.0640 0.0000 95.2640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.0640 0.0000 95.2640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.0640 0.0000 95.2640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.0640 0.0000 95.2640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[27]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[29]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.5920 0.0000 89.7920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.5920 0.0000 89.7920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.5920 0.0000 89.7920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.5920 0.0000 89.7920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.5920 0.0000 89.7920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[22]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 55.2650 131.4060 55.4650 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 55.2650 131.4060 55.4650 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 55.2650 131.4060 55.4650 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 55.2650 131.4060 55.4650 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 55.2650 131.4060 55.4650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.030936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.030936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.96053 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.10063 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 38.24046 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[0]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 9.8990 131.4060 10.0990 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 9.8990 131.4060 10.0990 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 9.8990 131.4060 10.0990 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 9.8990 131.4060 10.0990 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 9.8990 131.4060 10.0990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56742 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56742 LAYER M2 ;
    ANTENNAMAXAREACAR 11.76674 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.80361 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.84041 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.87714 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9110 0.2000 17.1110 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.9110 0.2000 17.1110 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.9110 0.2000 17.1110 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9110 0.2000 17.1110 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.9110 0.2000 17.1110 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.40684 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40684 LAYER M4 ;
    ANTENNAMAXAREACAR 13.07637 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.21759 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4450 0.2000 17.6450 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4450 0.2000 17.6450 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4450 0.2000 17.6450 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4450 0.2000 17.6450 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4450 0.2000 17.6450 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30916 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30916 LAYER M4 ;
    ANTENNAMAXAREACAR 12.51665 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 16.94857 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8980 0.2000 10.0980 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8980 0.2000 10.0980 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8980 0.2000 10.0980 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8980 0.2000 10.0980 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8980 0.2000 10.0980 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56742 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56742 LAYER M2 ;
    ANTENNAMAXAREACAR 11.76674 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.80361 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.84041 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.87714 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 41.2140 0.2000 41.4140 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 41.2140 0.2000 41.4140 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 41.2140 0.2000 41.4140 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 41.2140 0.2000 41.4140 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 41.2140 0.2000 41.4140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.028486 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.028486 LAYER M4 ;
    ANTENNAMAXAREACAR 51.90297 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 59.11859 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 46.4460 0.2000 46.6460 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 46.4460 0.2000 46.6460 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 46.4460 0.2000 46.6460 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 46.4460 0.2000 46.6460 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 46.4460 0.2000 46.6460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.030936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.030936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.96053 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.10063 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 38.24046 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 55.2660 0.2000 55.4660 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 55.2660 0.2000 55.4660 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 55.2660 0.2000 55.4660 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 55.2660 0.2000 55.4660 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 55.2660 0.2000 55.4660 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.030936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.030936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.96053 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.10063 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 38.24046 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 48.0380 0.2000 48.2380 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 48.0380 0.2000 48.2380 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 48.0380 0.2000 48.2380 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 48.0380 0.2000 48.2380 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 48.0380 0.2000 48.2380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.030936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.030936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.96053 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.10063 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 38.24046 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.2720 0.0000 103.4720 0.2000 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.3760 0.0000 107.5760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.3760 0.0000 107.5760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.3760 0.0000 107.5760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[16]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.7440 0.0000 108.9440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.7440 0.0000 108.9440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.7440 0.0000 108.9440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.7440 0.0000 108.9440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.7440 0.0000 108.9440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[8]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.1120 0.0000 110.3120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.1120 0.0000 110.3120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.1120 0.0000 110.3120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.1120 0.0000 110.3120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.1120 0.0000 110.3120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 41.2230 131.4060 41.4230 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 41.2230 131.4060 41.4230 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 41.2230 131.4060 41.4230 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 41.2230 131.4060 41.4230 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 41.2230 131.4060 41.4230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.064046 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.064046 LAYER M4 ;
    ANTENNAMAXAREACAR 53.5963 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 60.81181 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 46.4440 131.4060 46.6440 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 46.4440 131.4060 46.6440 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 46.4440 131.4060 46.6440 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 46.4440 131.4060 46.6440 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 46.4440 131.4060 46.6440 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.030936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.030936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.96053 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.10063 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 38.24046 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 48.0370 131.4060 48.2370 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 48.0370 131.4060 48.2370 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 48.0370 131.4060 48.2370 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 48.0370 131.4060 48.2370 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 48.0370 131.4060 48.2370 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.030936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.030936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.96053 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.10063 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 38.24046 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[1]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 17.3640 131.4060 17.5640 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 17.3640 131.4060 17.5640 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 17.3640 131.4060 17.5640 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 17.3640 131.4060 17.5640 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 17.3640 131.4060 17.5640 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.29968 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.29968 LAYER M4 ;
    ANTENNAMAXAREACAR 12.56501 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 16.99693 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 61.1440 0.2000 61.3440 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 61.1440 0.2000 61.3440 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 61.1440 0.2000 61.3440 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 61.1440 0.2000 61.3440 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 61.1440 0.2000 61.3440 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.235015 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.235015 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.938872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.938872 LAYER M2 ;
    ANTENNAMAXAREACAR 20.81647 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 28.31647 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.35878 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.40089 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 61.1460 131.4060 61.3460 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 61.1460 131.4060 61.3460 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 61.1460 131.4060 61.3460 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 61.1460 131.4060 61.3460 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 61.1460 131.4060 61.3460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.225565 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.225565 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.938872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.938872 LAYER M2 ;
    ANTENNAMAXAREACAR 20.81647 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 28.05829 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.10062 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.14274 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 16.9050 131.4060 17.1050 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 16.9050 131.4060 17.1050 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 16.9050 131.4060 17.1050 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 16.9050 131.4060 17.1050 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 16.9050 131.4060 17.1050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.424789 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.424789 LAYER M4 ;
    ANTENNAMAXAREACAR 13.53055 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.67173 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 2.8080 67.7440 3.1090 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9090 67.7440 2.2080 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.1090 67.7440 18.4090 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.8080 67.7440 57.1070 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.7080 67.7440 58.0070 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.6090 67.7440 58.9080 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.4080 67.7440 60.7070 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.7030 67.7440 130.0020 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.5090 67.7440 59.8090 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.8040 67.7440 129.1040 68.0440 ;
    END
    ANTENNADIFFAREA 108.1162 LAYER M5 ;
    ANTENNADIFFAREA 108.1162 LAYER M6 ;
    ANTENNADIFFAREA 108.1162 LAYER M7 ;
    ANTENNADIFFAREA 108.1162 LAYER M8 ;
    ANTENNADIFFAREA 108.1162 LAYER M9 ;
    ANTENNADIFFAREA 108.1162 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 120.6645 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 120.6645 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 784.3105 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 784.3105 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.1580 67.7440 4.4590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2580 67.7440 3.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3590 67.7440 2.6590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4580 67.7440 1.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0580 67.7440 5.3590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5580 67.7440 9.8590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6580 67.7440 8.9590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7590 67.7440 8.0580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8590 67.7440 7.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9590 67.7440 6.2590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3590 67.7440 11.6580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4590 67.7440 10.7590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0580 67.7440 14.3580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1590 67.7440 13.4590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2580 67.7440 12.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5580 67.7440 18.8590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6580 67.7440 17.9590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7580 67.7440 17.0590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8580 67.7440 16.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9590 67.7440 15.2580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2580 67.7440 21.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3590 67.7440 20.6590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1580 67.7440 22.4590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9590 67.7440 24.2580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0590 67.7440 23.3590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4590 67.7440 19.7590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7580 67.7440 26.0580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6590 67.7440 26.9590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5580 67.7440 27.8580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4590 67.7440 28.7590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8580 67.7440 25.1590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9590 67.7440 33.2590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1580 67.7440 31.4590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3590 67.7440 29.6580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2590 67.7440 30.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0580 67.7440 32.3590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8590 67.7440 34.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4580 67.7440 37.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6580 67.7440 35.9590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5580 67.7440 36.8590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3580 67.7440 38.6580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7590 67.7440 35.0580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8580 67.7440 43.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2590 67.7440 39.5590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1580 67.7440 40.4570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9580 67.7440 42.2580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0590 67.7440 41.3600 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3580 67.7440 47.6580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2590 67.7440 48.5590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4580 67.7440 46.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7590 67.7440 44.0590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5590 67.7440 45.8600 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6580 67.7440 44.9570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8580 67.7440 52.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1580 67.7440 49.4570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0590 67.7440 50.3600 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7590 67.7440 53.0590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9580 67.7440 51.2580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4580 67.7440 55.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5580 67.7440 54.8580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6580 67.7440 53.9580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3590 67.7440 56.6590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6570 67.7440 62.9570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7580 67.7440 62.0580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8580 67.7440 61.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1570 67.7440 67.4570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2580 67.7440 66.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3570 67.7440 65.6570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4570 67.7440 64.7570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5580 67.7440 63.8580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6580 67.7440 71.9580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7590 67.7440 71.0590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8570 67.7440 70.1570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9570 67.7440 69.2570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0580 67.7440 68.3580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1570 67.7440 76.4570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2580 67.7440 75.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3580 67.7440 74.6580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4580 67.7440 73.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.0580 67.7440 77.3580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5590 67.7440 72.8590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6580 67.7440 80.9580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7590 67.7440 80.0590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8570 67.7440 79.1570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9570 67.7440 78.2570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5590 67.7440 81.8590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.9570 67.7440 87.2570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1570 67.7440 85.4570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2580 67.7440 84.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3580 67.7440 83.6580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4580 67.7440 82.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0580 67.7440 86.3580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.4580 67.7440 91.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.5580 67.7440 90.8580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.6580 67.7440 89.9580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.8580 67.7440 88.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.7590 67.7440 89.0590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.0580 67.7440 95.3580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.1570 67.7440 94.4570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.3570 67.7440 92.6570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.9590 67.7440 96.2590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.2580 67.7440 93.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.3570 67.7440 101.6570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.5570 67.7440 99.8570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.6580 67.7440 98.9580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.7580 67.7440 98.0580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.8580 67.7440 97.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.4580 67.7440 100.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.8590 67.7440 106.1590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.9590 67.7440 105.2590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.0590 67.7440 104.3590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.2590 67.7440 102.5590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.1600 67.7440 103.4600 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.4580 67.7440 109.7580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.5580 67.7440 108.8580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.7580 67.7440 107.0580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.3590 67.7440 110.6590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.6590 67.7440 107.9590 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.9570 67.7440 114.2570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.0580 67.7440 113.3580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.1580 67.7440 112.4580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.2580 67.7440 111.5580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.8580 67.7440 115.1580 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.7570 67.7440 116.0570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.5570 67.7440 117.8570 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.2560 67.7440 120.5560 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.3560 67.7440 119.6560 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.4560 67.7440 118.7560 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.6560 67.7440 116.9560 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.7550 67.7440 125.0550 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.0560 67.7440 122.3560 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.8540 67.7440 124.1540 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.9550 67.7440 123.2550 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.6540 67.7440 125.9540 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.5540 67.7440 126.8540 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.4540 67.7440 127.7540 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.3530 67.7440 128.6530 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.1530 67.7440 130.4530 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.2540 67.7440 129.5540 68.0440 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.1550 67.7440 121.4550 68.0440 ;
    END
    ANTENNADIFFAREA 396.4798 LAYER M5 ;
    ANTENNADIFFAREA 396.4798 LAYER M6 ;
    ANTENNADIFFAREA 396.4798 LAYER M7 ;
    ANTENNADIFFAREA 396.4798 LAYER M8 ;
    ANTENNADIFFAREA 396.4798 LAYER M9 ;
    ANTENNADIFFAREA 396.4798 LAYER MRDL ;
    ANTENNAGATEAREA 40.353 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 3726.063 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3726.063 LAYER M5 ;
    ANTENNAMAXAREACAR 175.1118 LAYER M5 ;
    ANTENNAGATEAREA 40.353 LAYER M6 ;
    ANTENNAGATEAREA 40.353 LAYER M7 ;
    ANTENNAGATEAREA 40.353 LAYER M8 ;
    ANTENNAGATEAREA 40.353 LAYER M9 ;
    ANTENNAGATEAREA 40.353 LAYER MRDL ;
  END VSS

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.3760 0.0000 107.5760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.3760 0.0000 107.5760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[16]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 103.2720 0.0000 103.4720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.2720 0.0000 103.4720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.2720 0.0000 103.4720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.2720 0.0000 103.4720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[10]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[19]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8940 0.0000 25.0940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8940 0.0000 25.0940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8940 0.0000 25.0940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8940 0.0000 25.0940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8940 0.0000 25.0940 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[30]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2630 0.0000 26.4630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2630 0.0000 26.4630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2630 0.0000 26.4630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2630 0.0000 26.4630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2630 0.0000 26.4630 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 57.9930 0.2000 58.1930 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 57.9930 0.2000 58.1930 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 57.9930 0.2000 58.1930 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 57.9930 0.2000 58.1930 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 57.9930 0.2000 58.1930 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16336 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16336 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.244428 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.244428 LAYER M2 ;
    ANTENNAMAXAREACAR 12.92088 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.195923 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.195923 LAYER M3 ;
    ANTENNAMAXAREACAR 27.54596 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 42.46913 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 45.79089 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.5178 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.8762 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8762 LAYER M2 ;
    ANTENNAMAXAREACAR 6.520677 LAYER M2 ;
    ANTENNAGATEAREA 0.5178 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 6.813024 LAYER M3 ;
    ANTENNAGATEAREA 0.5178 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.105351 LAYER M4 ;
    ANTENNAGATEAREA 0.5178 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.39766 LAYER M5 ;
    ANTENNAGATEAREA 0.5178 LAYER M6 ;
    ANTENNAGATEAREA 0.5178 LAYER M7 ;
    ANTENNAGATEAREA 0.5178 LAYER M8 ;
    ANTENNAGATEAREA 0.5178 LAYER M9 ;
    ANTENNAGATEAREA 0.5178 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.5178 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.88202 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.88202 LAYER M2 ;
    ANTENNAMAXAREACAR 6.531917 LAYER M2 ;
    ANTENNAGATEAREA 0.5178 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 6.824263 LAYER M3 ;
    ANTENNAGATEAREA 0.5178 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.11659 LAYER M4 ;
    ANTENNAGATEAREA 0.5178 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.408897 LAYER M5 ;
    ANTENNAGATEAREA 0.5178 LAYER M6 ;
    ANTENNAGATEAREA 0.5178 LAYER M7 ;
    ANTENNAGATEAREA 0.5178 LAYER M8 ;
    ANTENNAGATEAREA 0.5178 LAYER M9 ;
    ANTENNAGATEAREA 0.5178 LAYER MRDL ;
  END OEB1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 57.6400 131.4060 57.8400 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 57.6400 131.4060 57.8400 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 57.6400 131.4060 57.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 57.6400 131.4060 57.8400 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 57.6400 131.4060 57.8400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.269868 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.269868 LAYER M2 ;
    ANTENNAMAXAREACAR 14.18107 LAYER M2 ;
    ANTENNAGATEAREA 0.0792 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 7.855984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.855984 LAYER M3 ;
    ANTENNAMAXAREACAR 102.1479 LAYER M3 ;
    ANTENNAGATEAREA 0.0792 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 115.2794 LAYER M4 ;
    ANTENNAGATEAREA 0.0792 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 117.186 LAYER M5 ;
    ANTENNAGATEAREA 0.0792 LAYER M6 ;
    ANTENNAGATEAREA 0.0792 LAYER M7 ;
    ANTENNAGATEAREA 0.0792 LAYER M8 ;
    ANTENNAGATEAREA 0.0792 LAYER M9 ;
    ANTENNAGATEAREA 0.0792 LAYER MRDL ;
  END SD

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.3100 0.0000 41.5100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.3100 0.0000 41.5100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.3100 0.0000 41.5100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.3100 0.0000 41.5100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.3100 0.0000 41.5100 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9420 0.0000 40.1420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9420 0.0000 40.1420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9420 0.0000 40.1420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9420 0.0000 40.1420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9420 0.0000 40.1420 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[23]

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 57.9830 131.4060 58.1830 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 57.9830 131.4060 58.1830 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 57.9830 131.4060 58.1830 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 57.9830 131.4060 58.1830 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 57.9830 131.4060 58.1830 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.236068 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.236068 LAYER M2 ;
    ANTENNAMAXAREACAR 12.52839 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 7.521058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.521058 LAYER M3 ;
    ANTENNAMAXAREACAR 166.5476 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 180.7327 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 184.0013 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS1

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8120 0.0000 34.0120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8120 0.0000 34.0120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8120 0.0000 34.0120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8120 0.0000 34.0120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8120 0.0000 34.0120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[28]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 0.0000 33.3020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 0.0000 33.3020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 0.0000 33.3020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 0.0000 33.3020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 0.0000 33.3020 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.2050 0.0000 37.4050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.2050 0.0000 37.4050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.2050 0.0000 37.4050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.2050 0.0000 37.4050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.2050 0.0000 37.4050 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[25]

  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4700 0.0000 34.6700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4700 0.0000 34.6700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4700 0.0000 34.6700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4700 0.0000 34.6700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4700 0.0000 34.6700 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[28]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8380 0.0000 36.0380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8380 0.0000 36.0380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8380 0.0000 36.0380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8380 0.0000 36.0380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8380 0.0000 36.0380 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[11]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6300 0.0000 27.8300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6300 0.0000 27.8300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6300 0.0000 27.8300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6300 0.0000 27.8300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6300 0.0000 27.8300 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[19]

  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9980 0.0000 29.1980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9980 0.0000 29.1980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9980 0.0000 29.1980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9980 0.0000 29.1980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9980 0.0000 29.1980 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[30]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3660 0.0000 30.5660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3660 0.0000 30.5660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3660 0.0000 30.5660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3660 0.0000 30.5660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3660 0.0000 30.5660 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7340 0.0000 31.9340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7340 0.0000 31.9340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7340 0.0000 31.9340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7340 0.0000 31.9340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7340 0.0000 31.9340 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.5360 0.0000 100.7360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.5360 0.0000 100.7360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.5360 0.0000 100.7360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.5360 0.0000 100.7360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.5360 0.0000 100.7360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[18]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[31]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[20]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[24]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[27]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.5180 0.0000 49.7180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.5180 0.0000 49.7180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.5180 0.0000 49.7180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.5180 0.0000 49.7180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.5180 0.0000 49.7180 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[15]

  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8860 0.0000 51.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8860 0.0000 51.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8860 0.0000 51.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8860 0.0000 51.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8860 0.0000 51.0860 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[27]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[21]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[15]

  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7830 0.0000 46.9830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7830 0.0000 46.9830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7830 0.0000 46.9830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7830 0.0000 46.9830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7830 0.0000 46.9830 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[29]

  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1500 0.0000 48.3500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1500 0.0000 48.3500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1500 0.0000 48.3500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1500 0.0000 48.3500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1500 0.0000 48.3500 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[21]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[29]

  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.4140 0.0000 45.6140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.4140 0.0000 45.6140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.4140 0.0000 45.6140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.4140 0.0000 45.6140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.4140 0.0000 45.6140 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[22]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[26]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[22]

  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6780 0.0000 42.8780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6780 0.0000 42.8780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6780 0.0000 42.8780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6780 0.0000 42.8780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6780 0.0000 42.8780 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[31]

  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0460 0.0000 44.2460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0460 0.0000 44.2460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0460 0.0000 44.2460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0460 0.0000 44.2460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0460 0.0000 44.2460 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[26]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[23]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5740 0.0000 38.7740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5740 0.0000 38.7740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5740 0.0000 38.7740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5740 0.0000 38.7740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5740 0.0000 38.7740 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[25]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.4140 -0.0020 68.6140 0.1980 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.4140 -0.0020 68.6140 0.1980 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.4140 -0.0020 68.6140 0.1980 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.4140 -0.0020 68.6140 0.1980 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.4140 -0.0020 68.6140 0.1980 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28848 LAYER M3 ;
    ANTENNAMAXAREACAR 62.60445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81937 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.03381 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[16]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.8300 0.0000 62.0300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.8300 0.0000 62.0300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.8300 0.0000 62.0300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.8300 0.0000 62.0300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.8300 0.0000 62.0300 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1980 0.0000 63.3980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1980 0.0000 63.3980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1980 0.0000 63.3980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1980 0.0000 63.3980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1980 0.0000 63.3980 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[16]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5660 0.0000 64.7660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5660 0.0000 64.7660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5660 0.0000 64.7660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5660 0.0000 64.7660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5660 0.0000 64.7660 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[17]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0940 0.0000 59.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0940 0.0000 59.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0940 0.0000 59.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0940 0.0000 59.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0940 0.0000 59.2940 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4620 0.0000 60.6620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4620 0.0000 60.6620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4620 0.0000 60.6620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4620 0.0000 60.6620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4620 0.0000 60.6620 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3580 0.0000 56.5580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3580 0.0000 56.5580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3580 0.0000 56.5580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3580 0.0000 56.5580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3580 0.0000 56.5580 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[18]

  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.7260 0.0000 57.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.7260 0.0000 57.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.7260 0.0000 57.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.7260 0.0000 57.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.7260 0.0000 57.9260 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[17]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[18]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9900 0.0000 55.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9900 0.0000 55.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9900 0.0000 55.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9900 0.0000 55.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9900 0.0000 55.1900 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2540 0.0000 52.4540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2540 0.0000 52.4540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2540 0.0000 52.4540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2540 0.0000 52.4540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2540 0.0000 52.4540 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[20]

  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.6220 0.0000 53.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.6220 0.0000 53.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.6220 0.0000 53.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.6220 0.0000 53.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.6220 0.0000 53.8220 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[24]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.6480 0.0000 78.8480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.6480 0.0000 78.8480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.6480 0.0000 78.8480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.6480 0.0000 78.8480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.6480 0.0000 78.8480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[28]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.0160 0.0000 80.2160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.0160 0.0000 80.2160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.0160 0.0000 80.2160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.0160 0.0000 80.2160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.0160 0.0000 80.2160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[23]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.7520 0.0000 82.9520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.7520 0.0000 82.9520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.7520 0.0000 82.9520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.7520 0.0000 82.9520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.7520 0.0000 82.9520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[25]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[25]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.3840 0.0000 81.5840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.3840 0.0000 81.5840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.3840 0.0000 81.5840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.3840 0.0000 81.5840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.3840 0.0000 81.5840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28836 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28836 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.81366 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.0281 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[19]
  OBS
    LAYER M1 ;
      RECT 0.8000 42.0230 130.6060 47.4370 ;
      RECT 0.8000 42.0230 130.6060 47.4370 ;
      RECT 0.8000 42.0230 130.6060 47.4370 ;
      RECT 21.3780 0.0000 22.2680 0.8000 ;
      RECT 0.0000 58.7930 1.5010 60.5440 ;
      RECT 129.9050 58.7830 131.4060 60.5460 ;
      RECT 0.0000 56.0660 0.8000 57.3930 ;
      RECT 0.0000 45.8440 3.0010 45.8460 ;
      RECT 0.0000 61.9440 3.0010 61.9460 ;
      RECT 0.0000 54.6650 3.0010 54.6660 ;
      RECT 0.0000 47.2460 0.8000 47.4380 ;
      RECT 130.6060 56.0650 131.4060 57.0400 ;
      RECT 0.8000 48.8370 131.4060 51.8380 ;
      RECT 130.6060 47.2440 131.4060 47.4370 ;
      RECT 0.0000 10.6990 131.4060 16.3050 ;
      RECT 0.8000 40.6230 130.6060 42.0140 ;
      RECT 0.0000 16.3050 130.6060 16.3110 ;
      RECT 0.0000 10.6990 130.6060 16.3110 ;
      RECT 0.0000 10.6990 130.6060 16.3110 ;
      RECT 0.0000 10.6990 130.6060 16.3110 ;
      RECT 0.0000 18.2450 131.4060 40.6140 ;
      RECT 0.8000 40.6140 131.4060 40.6230 ;
      RECT 0.8000 18.2450 131.4060 40.6230 ;
      RECT 0.8000 18.2450 131.4060 40.6230 ;
      RECT 0.8000 18.2450 131.4060 40.6230 ;
      RECT 0.8000 18.1640 131.4060 40.6140 ;
      RECT 0.8000 18.1640 131.4060 40.6140 ;
      RECT 0.8000 18.1640 131.4060 40.6140 ;
      RECT 0.8000 16.3110 130.6060 40.6140 ;
      RECT 0.8000 16.3110 130.6060 40.6140 ;
      RECT 0.8000 16.3110 130.6060 40.6140 ;
      RECT 0.8000 18.1640 131.4060 18.2450 ;
      RECT 0.8000 16.3110 130.6060 18.1640 ;
      RECT 0.0000 10.6980 130.6060 16.3050 ;
      RECT 0.0000 10.6980 130.6060 16.3050 ;
      RECT 0.0000 10.6980 130.6060 16.3050 ;
      RECT 0.0000 10.6980 130.6060 10.6990 ;
      RECT 0.0000 0.0000 19.9780 9.2980 ;
      RECT 0.0000 0.0000 19.9780 0.8000 ;
      RECT 0.8000 9.2990 130.6060 10.6980 ;
      RECT 0.8000 9.2980 131.4060 9.2990 ;
      RECT 0.0000 0.8000 131.4060 9.2980 ;
      RECT 0.8000 0.8000 130.6060 10.6980 ;
      RECT 0.8000 0.8000 130.6060 10.6980 ;
      RECT 0.8000 0.8000 130.6060 10.6980 ;
      RECT 0.8000 0.8000 131.4060 9.2990 ;
      RECT 0.8000 0.8000 131.4060 9.2990 ;
      RECT 0.8000 0.8000 131.4060 9.2990 ;
      RECT 111.4180 0.0000 131.4060 9.2980 ;
      RECT 111.4180 0.0000 131.4060 0.8000 ;
      RECT 0.0000 42.0230 131.4060 45.8440 ;
      RECT 0.0000 42.0140 130.6060 45.8440 ;
      RECT 0.0000 42.0140 130.6060 45.8440 ;
      RECT 0.0000 42.0140 130.6060 45.8440 ;
      RECT 0.0000 42.0140 130.6060 42.0230 ;
      RECT 0.0000 61.9460 131.4060 68.0440 ;
      RECT 0.8000 58.7930 130.6060 61.9460 ;
      RECT 0.8000 57.3930 130.6060 61.9460 ;
      RECT 0.8000 57.3930 130.6060 60.5460 ;
      RECT 0.8000 57.3930 130.6060 60.5460 ;
      RECT 0.8000 57.3930 130.6060 60.5460 ;
      RECT 0.8000 57.3930 130.6060 60.5460 ;
      RECT 0.8000 57.3930 130.6060 60.5460 ;
      RECT 0.8000 57.3930 130.6060 60.5440 ;
      RECT 0.8000 57.3930 130.6060 60.5440 ;
      RECT 0.8000 57.3930 130.6060 60.5440 ;
      RECT 0.8000 57.3930 130.6060 60.5440 ;
      RECT 0.8000 57.3930 130.6060 60.5440 ;
      RECT 0.8000 54.6660 130.6060 61.9440 ;
      RECT 0.8000 54.6660 130.6060 61.9440 ;
      RECT 0.8000 54.6660 130.6060 60.5460 ;
      RECT 0.8000 54.6660 130.6060 60.5460 ;
      RECT 0.8000 54.6660 130.6060 60.5460 ;
      RECT 0.8000 54.6660 130.6060 60.5460 ;
      RECT 0.8000 54.6660 130.6060 60.5440 ;
      RECT 0.8000 57.0400 130.6060 57.3930 ;
      RECT 0.0000 48.8380 131.4060 54.6650 ;
      RECT 0.8000 48.8380 130.6060 61.9440 ;
      RECT 0.8000 48.8380 130.6060 61.9440 ;
      RECT 0.8000 48.8380 130.6060 60.5460 ;
      RECT 0.8000 48.8380 130.6060 60.5460 ;
      RECT 0.8000 48.8380 130.6060 60.5440 ;
      RECT 0.8000 48.8380 130.6060 60.5440 ;
      RECT 0.8000 48.8380 130.6060 60.5440 ;
      RECT 0.8000 48.8380 130.6060 60.5440 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 48.8380 130.6060 57.3930 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 48.8370 ;
      RECT 0.8000 42.0230 130.6060 47.4370 ;
      RECT 0.8000 42.0230 130.6060 47.4370 ;
    LAYER PO ;
      RECT 0.0000 0.0000 131.4060 68.0440 ;
    LAYER M2 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8830 ;
      RECT 0.9000 48.9380 130.5060 58.8830 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 58.8930 1.5010 60.4440 ;
      RECT 0.0000 56.1660 0.9000 57.2930 ;
      RECT 0.0000 54.5650 3.0010 54.5660 ;
      RECT 0.0000 62.0440 3.0010 62.0460 ;
      RECT 130.5060 56.1650 131.4060 56.9400 ;
      RECT 129.9050 58.8830 131.4060 60.4460 ;
      RECT 0.9000 45.7460 130.5060 48.9370 ;
      RECT 0.0000 0.0000 19.8780 9.1980 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 45.7440 130.5060 45.7460 ;
      RECT 0.0000 42.1230 130.5060 45.7460 ;
      RECT 0.0000 42.1230 131.4060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 42.1230 ;
      RECT 0.9000 42.1230 130.5060 48.9370 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 42.1140 ;
      RECT 0.0000 18.3450 131.4060 40.5140 ;
      RECT 0.9000 40.5140 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 18.3450 ;
      RECT 0.9000 16.2110 130.5060 18.2640 ;
      RECT 0.0000 16.2050 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 131.4060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 10.7990 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 10.7980 ;
      RECT 0.9000 9.1980 131.4060 9.1990 ;
      RECT 0.0000 0.9000 131.4060 9.1980 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 111.5180 0.0000 131.4060 9.1980 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 48.9380 131.4060 54.5650 ;
      RECT 0.9000 48.9370 131.4060 48.9380 ;
      RECT 0.9000 45.7460 130.5060 48.9380 ;
      RECT 0.0000 62.0460 131.4060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 54.5660 130.5060 60.4460 ;
      RECT 0.9000 48.9380 130.5060 60.4460 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
    LAYER M3 ;
      RECT 0.9000 45.7460 130.5060 48.9380 ;
      RECT 0.0000 62.0460 131.4060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 54.5660 130.5060 60.4460 ;
      RECT 0.9000 48.9380 130.5060 60.4460 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8830 ;
      RECT 0.9000 48.9380 130.5060 58.8830 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 62.0440 3.0010 62.0460 ;
      RECT 0.0000 54.5650 3.0010 54.5660 ;
      RECT 0.0000 56.1660 0.9000 57.2930 ;
      RECT 0.0000 58.8930 1.5010 60.4440 ;
      RECT 129.9050 58.8830 131.4060 60.4460 ;
      RECT 130.5060 56.1650 131.4060 56.9400 ;
      RECT 0.9000 45.7460 130.5060 48.9370 ;
      RECT 0.0000 0.0000 19.8780 9.1980 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 45.7440 130.5060 45.7460 ;
      RECT 0.0000 42.1230 130.5060 45.7460 ;
      RECT 0.0000 42.1230 131.4060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 42.1230 ;
      RECT 0.9000 42.1230 130.5060 48.9370 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 42.1140 ;
      RECT 0.0000 18.3450 131.4060 40.5140 ;
      RECT 0.9000 40.5140 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 18.3450 ;
      RECT 0.9000 16.2110 130.5060 18.2640 ;
      RECT 0.0000 16.2050 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 131.4060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 10.7990 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 10.7980 ;
      RECT 0.9000 9.1980 131.4060 9.1990 ;
      RECT 0.0000 0.9000 131.4060 9.1980 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 111.5180 0.0000 131.4060 9.1980 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 48.9380 131.4060 54.5650 ;
      RECT 0.9000 48.9370 131.4060 48.9380 ;
    LAYER M4 ;
      RECT 0.0000 16.2050 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 131.4060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 10.7990 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 16.2050 ;
      RECT 0.9000 9.1990 130.5060 10.7980 ;
      RECT 0.9000 9.1980 131.4060 9.1990 ;
      RECT 0.0000 0.9000 131.4060 9.1980 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 111.5180 0.0000 131.4060 9.1980 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 48.9380 131.4060 54.5650 ;
      RECT 0.9000 48.9370 131.4060 48.9380 ;
      RECT 0.9000 45.7460 130.5060 48.9380 ;
      RECT 0.0000 62.0460 131.4060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 68.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 54.5660 130.5060 60.4460 ;
      RECT 0.9000 48.9380 130.5060 60.4460 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 48.9380 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8930 ;
      RECT 0.9000 48.9380 130.5060 58.8830 ;
      RECT 0.9000 48.9380 130.5060 58.8830 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 62.0440 3.0010 62.0460 ;
      RECT 0.0000 54.5650 3.0010 54.5660 ;
      RECT 0.0000 56.1660 0.9000 57.2930 ;
      RECT 0.0000 58.8930 1.5010 60.4440 ;
      RECT 129.9050 58.8830 131.4060 60.4460 ;
      RECT 130.5060 56.1650 131.4060 56.9400 ;
      RECT 0.9000 45.7460 130.5060 48.9370 ;
      RECT 0.0000 0.0000 19.8780 9.1980 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 45.7440 130.5060 45.7460 ;
      RECT 0.0000 42.1230 130.5060 45.7460 ;
      RECT 0.0000 42.1230 131.4060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 42.1230 ;
      RECT 0.9000 42.1230 130.5060 48.9370 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 45.7440 ;
      RECT 0.9000 40.5230 130.5060 42.1140 ;
      RECT 0.0000 18.3450 131.4060 40.5140 ;
      RECT 0.9000 40.5140 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 18.3450 ;
      RECT 0.9000 16.2110 130.5060 18.2640 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 131.4060 68.0440 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 131.4060 68.0440 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 131.4060 68.0440 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 131.4060 68.0440 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 131.4060 68.0440 ;
    LAYER M5 ;
      RECT 131.1530 67.0440 131.4060 68.0440 ;
      RECT 0.0000 67.0440 0.7580 68.0440 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 62.0440 3.0010 62.0460 ;
      RECT 0.0000 56.1660 0.9000 57.2930 ;
      RECT 0.0000 51.5650 130.5060 54.5660 ;
      RECT 0.0000 58.8930 1.5010 60.4440 ;
      RECT 129.9050 58.8830 131.4060 60.4460 ;
      RECT 130.5060 56.1650 131.4060 56.9400 ;
      RECT 0.0000 10.7990 131.4060 16.2050 ;
      RECT 0.0000 42.1230 131.4060 45.7440 ;
      RECT 0.0000 45.7440 130.5060 45.7460 ;
      RECT 0.0000 42.1230 130.5060 45.7460 ;
      RECT 0.9000 45.7460 130.5060 48.9370 ;
      RECT 0.9000 42.1230 130.5060 48.9370 ;
      RECT 0.0000 16.2050 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.0000 10.7990 130.5060 16.2110 ;
      RECT 0.9000 16.2110 130.5060 18.2640 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 45.7440 ;
      RECT 0.0000 42.1140 130.5060 42.1230 ;
      RECT 0.0000 18.3450 131.4060 40.5140 ;
      RECT 0.9000 40.5230 130.5060 42.1140 ;
      RECT 0.9000 18.3450 130.5060 42.1140 ;
      RECT 0.9000 18.3450 130.5060 42.1140 ;
      RECT 0.9000 18.3450 130.5060 42.1140 ;
      RECT 0.9000 40.5140 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.3450 131.4060 40.5230 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 16.2110 130.5060 40.5140 ;
      RECT 0.9000 18.2640 131.4060 18.3450 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 16.2050 ;
      RECT 0.0000 10.7980 130.5060 10.7990 ;
      RECT 0.0000 0.0000 19.8780 9.1980 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.9000 9.1990 130.5060 10.7980 ;
      RECT 0.0000 0.9000 131.4060 9.1980 ;
      RECT 0.9000 0.9000 130.5060 10.7980 ;
      RECT 0.9000 0.9000 130.5060 10.7980 ;
      RECT 0.9000 0.9000 130.5060 10.7980 ;
      RECT 0.9000 9.1980 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 0.9000 0.9000 131.4060 9.1990 ;
      RECT 111.5180 0.0000 131.4060 9.1980 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 62.0460 131.4060 67.0440 ;
      RECT 0.0000 48.9380 131.4060 54.5650 ;
      RECT 0.9000 48.9370 131.4060 48.9380 ;
      RECT 0.9000 45.7460 130.5060 48.9380 ;
      RECT 0.9000 58.8930 130.5060 62.0460 ;
      RECT 0.9000 57.2930 130.5060 62.0460 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 58.8930 130.5060 62.0440 ;
      RECT 0.9000 57.2930 130.5060 60.4460 ;
      RECT 0.9000 57.2930 130.5060 60.4460 ;
      RECT 0.9000 57.2930 130.5060 60.4460 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 57.2930 130.5060 60.4440 ;
      RECT 0.9000 56.1650 130.5060 60.4460 ;
      RECT 0.9000 56.1650 130.5060 60.4460 ;
      RECT 0.9000 56.1650 130.5060 60.4440 ;
      RECT 0.9000 56.1650 130.5060 60.4440 ;
      RECT 0.9000 56.1650 130.5060 60.4440 ;
      RECT 0.9000 56.1650 130.5060 60.4440 ;
      RECT 0.9000 56.1650 130.5060 60.4440 ;
      RECT 0.9000 56.1650 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 60.4440 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8930 ;
      RECT 0.9000 54.5660 130.5060 58.8830 ;
      RECT 0.9000 56.9400 130.5060 57.2930 ;
  END
END SRAMLP2RW16x32

MACRO unitTile
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0 BY 0 ;
  SYMMETRY X Y R90 ;
END unitTile

MACRO SRAMLP2RW32x4
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 55.645 BY 64.819 ;
  SYMMETRY X Y R90 ;

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 40.0630 0.2000 40.2630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 25.1380 55.6450 25.3380 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 25.1380 55.6450 25.3380 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 25.1380 55.6450 25.3380 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 25.1380 55.6450 25.3380 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 25.1380 55.6450 25.3380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 32.7080 55.6450 32.9080 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 31.2190 55.6450 31.4190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 40.0490 55.6450 40.2490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 16.7920 55.6450 16.9920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 17.2990 55.6450 17.4990 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 17.2990 55.6450 17.4990 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 17.2990 55.6450 17.4990 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 17.2990 55.6450 17.4990 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 17.2990 55.6450 17.4990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE1

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 25.9140 55.6450 26.1140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.0260 0.0000 34.2260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O1[1]

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.1070 0.0000 21.3070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 9.7790 55.6450 9.9790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB1

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 30.5900 0.2000 30.7900 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 30.5900 0.2000 30.7900 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 30.5900 0.2000 30.7900 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 30.5900 0.2000 30.7900 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 30.5900 0.2000 30.7900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.5160 64.5190 10.8170 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.4160 64.5190 11.7170 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.1160 64.5190 23.4150 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.0150 64.5190 24.3140 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.6140 64.5190 45.9150 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.5160 64.5190 46.8160 64.8190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.5390 0.0000 34.7390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.7800 0.2000 9.9800 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.9160 64.5190 7.2150 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.8160 64.5190 8.1150 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.8170 64.5190 17.1160 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.7170 64.5190 18.0170 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.3170 64.5190 48.6170 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.2170 64.5190 49.5160 64.8190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDD

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.8020 0.0000 27.0020 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.191048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191048 LAYER M3 ;
  END O2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.4990 0.0000 27.6990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.7630 0.0000 24.9630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[2]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.1310 0.0000 26.3310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[0]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.6370 0.0000 30.8370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[2]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.5720 0.0000 28.7720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 39.02243 LAYER M4 ;
    ANTENNADIFFAREA 39.02243 LAYER M5 ;
    ANTENNADIFFAREA 39.02243 LAYER M6 ;
    ANTENNADIFFAREA 39.02243 LAYER M7 ;
    ANTENNADIFFAREA 39.02243 LAYER M8 ;
    ANTENNADIFFAREA 39.02243 LAYER M9 ;
    ANTENNADIFFAREA 39.02243 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.215168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.215168 LAYER M3 ;
    ANTENNAGATEAREA 4.887 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 83.50632 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 83.50632 LAYER M4 ;
    ANTENNAMAXAREACAR 60.60049 LAYER M4 ;
    ANTENNAGATEAREA 4.887 LAYER M5 ;
    ANTENNAGATEAREA 4.887 LAYER M6 ;
    ANTENNAGATEAREA 4.887 LAYER M7 ;
    ANTENNAGATEAREA 4.887 LAYER M8 ;
    ANTENNAGATEAREA 4.887 LAYER M9 ;
    ANTENNAGATEAREA 4.887 LAYER MRDL ;
  END O2[1]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.9400 0.0000 30.1400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.191048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191048 LAYER M3 ;
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.3080 0.0000 31.5080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.191048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191048 LAYER M3 ;
  END O1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.2690 0.0000 29.4690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[3]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.3730 0.0000 33.5730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.6760 0.0000 32.8760 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.0050 0.0000 32.2050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[0]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.2460 0.2000 17.4460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.7860 0.2000 16.9860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB2

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 32.7220 0.2000 32.9220 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 31.2330 0.2000 31.4330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 54.4290 55.6450 54.6290 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 54.4290 55.6450 54.6290 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 54.4290 55.6450 54.6290 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 54.4290 55.6450 54.6290 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 54.4290 55.6450 54.6290 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 57.9120 55.6450 58.1120 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 57.9120 55.6450 58.1120 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 57.9120 55.6450 58.1120 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 57.9120 55.6450 58.1120 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 57.9120 55.6450 58.1120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.4340 0.0000 25.6340 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.191048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191048 LAYER M3 ;
  END O2[2]

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 57.9590 0.2000 58.1590 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 57.9590 0.2000 58.1590 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 57.9590 0.2000 58.1590 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 57.9590 0.2000 58.1590 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 57.9590 0.2000 58.1590 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4450 54.7830 55.6450 54.9830 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4450 54.7830 55.6450 54.9830 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4450 54.7830 55.6450 54.9830 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4450 54.7830 55.6450 54.9830 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4450 54.7830 55.6450 54.9830 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS1

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 54.7690 0.2000 54.9690 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 54.7690 0.2000 54.9690 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 54.7690 0.2000 54.9690 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 54.7690 0.2000 54.9690 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 54.7690 0.2000 54.9690 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 25.9280 0.2000 26.1280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[4]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.3950 0.0000 23.5950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[3]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.0660 0.0000 24.2660 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.191048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191048 LAYER M3 ;
  END O2[3]

  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.3660 64.5190 16.6670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.0660 64.5190 46.3660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.7670 64.5190 13.0670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.1670 64.5190 45.4670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.5670 64.5190 14.8660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.9670 64.5190 47.2660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.4660 64.5190 15.7660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.6660 64.5190 13.9660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.2660 64.5190 44.5660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8660 64.5190 12.1660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.3670 64.5190 43.6660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.5660 64.5190 32.8650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.9670 64.5190 11.2660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.4670 64.5190 42.7670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.6660 64.5190 31.9660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.0670 64.5190 10.3670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.5660 64.5190 41.8670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.7650 64.5190 31.0660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.1660 64.5190 9.4670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.8670 64.5190 39.1660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.0660 64.5190 28.3650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.4670 64.5190 6.7660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.9670 64.5190 38.2670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.1660 64.5190 27.4660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.5670 64.5190 5.8670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.7670 64.5190 40.0660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.9660 64.5190 29.2650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.6660 64.5190 40.9670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.8650 64.5190 30.1660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.2660 64.5190 8.5670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.2660 64.5190 35.5660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.4650 64.5190 24.7650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.8660 64.5190 3.1660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.3670 64.5190 34.6670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.5660 64.5190 23.8660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9670 64.5190 2.2670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.4660 64.5190 33.7660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.6650 64.5190 22.9650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.0650 64.5190 1.3650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.0660 64.5190 37.3670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.2650 64.5190 26.5660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.6660 64.5190 4.9670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.1660 64.5190 36.4670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.3650 64.5190 25.6660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.7660 64.5190 4.0670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.1650 64.5190 54.4650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.7650 64.5190 22.0650 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.3670 64.5190 52.6670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.9670 64.5190 20.2670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.2660 64.5190 53.5660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.8660 64.5190 21.1660 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.4670 64.5190 51.7670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.0670 64.5190 19.3670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.5660 64.5190 50.8670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.1660 64.5190 18.4670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.6660 64.5190 49.9670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.2660 64.5190 17.5670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.7660 64.5190 49.0670 64.8190 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.8660 64.5190 48.1660 64.8190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0000 0.8000 54.8450 9.1800 ;
      RECT 0.0000 0.8000 54.8450 9.1800 ;
      RECT 0.0000 0.8000 55.6450 9.1790 ;
      RECT 0.8000 0.8000 54.8450 10.5790 ;
      RECT 0.8000 0.8000 54.8450 10.5790 ;
      RECT 0.8000 0.8000 54.8450 10.5790 ;
      RECT 35.3390 0.0000 55.6450 9.1790 ;
      RECT 35.3390 0.0000 55.6450 0.8000 ;
      RECT 0.0000 40.8630 55.6450 53.8290 ;
      RECT 0.8000 40.8490 55.6450 53.8290 ;
      RECT 0.8000 40.8490 55.6450 53.8290 ;
      RECT 0.8000 40.8490 55.6450 53.8290 ;
      RECT 0.8000 40.8490 55.6450 40.8630 ;
      RECT 0.8000 57.3120 54.8450 57.3590 ;
      RECT 0.0000 26.7280 55.6450 29.9900 ;
      RECT 0.8000 26.7280 54.8450 32.1080 ;
      RECT 0.8000 26.7280 54.8450 32.1080 ;
      RECT 0.8000 26.7280 54.8450 32.1080 ;
      RECT 0.8000 26.7280 54.8450 32.1080 ;
      RECT 0.8000 26.7280 54.8450 32.1080 ;
      RECT 0.8000 26.7280 54.8450 32.1080 ;
      RECT 0.8000 26.7140 55.6450 29.9900 ;
      RECT 0.8000 26.7140 55.6450 29.9900 ;
      RECT 0.8000 26.7140 55.6450 29.9900 ;
      RECT 0.8000 26.7140 55.6450 26.7280 ;
      RECT 0.8000 32.1080 54.8450 32.1220 ;
      RECT 0.8000 26.7280 54.8450 32.1220 ;
      RECT 0.8000 26.7280 54.8450 32.1220 ;
      RECT 0.8000 26.7280 54.8450 32.1220 ;
      RECT 0.8000 26.7280 54.8450 32.1220 ;
      RECT 0.8000 26.7280 54.8450 32.1220 ;
      RECT 0.8000 26.7280 54.8450 32.1220 ;
      RECT 0.0000 58.7590 55.6450 64.8190 ;
      RECT 0.8000 55.5690 54.8450 58.7120 ;
      RECT 0.8000 55.5690 54.8450 58.7120 ;
      RECT 0.8000 55.5690 54.8450 58.7120 ;
      RECT 0.8000 55.5690 54.8450 58.7120 ;
      RECT 0.8000 55.5830 54.8450 58.7120 ;
      RECT 0.8000 55.5690 54.8450 58.7120 ;
      RECT 0.8000 54.1690 54.8450 58.7120 ;
      RECT 0.8000 54.1690 54.8450 58.7120 ;
      RECT 0.8000 54.1690 54.8450 58.7120 ;
      RECT 0.8000 54.1690 54.8450 58.7120 ;
      RECT 0.8000 54.1690 54.8450 58.7120 ;
      RECT 0.0000 33.5220 54.8450 39.4630 ;
      RECT 0.0000 33.5220 54.8450 39.4630 ;
      RECT 0.0000 33.5220 54.8450 39.4630 ;
      RECT 0.0000 39.4490 54.8450 39.4630 ;
      RECT 0.0000 33.5220 55.6450 39.4490 ;
      RECT 0.8000 33.5220 54.8450 40.8490 ;
      RECT 0.8000 33.5220 54.8450 40.8490 ;
      RECT 0.8000 33.5220 54.8450 40.8490 ;
      RECT 21.9070 0.0000 22.7950 0.8000 ;
      RECT 54.1440 55.5830 55.6450 57.3120 ;
      RECT 0.0000 51.1680 54.8450 54.1690 ;
      RECT 52.6440 29.9900 55.6450 30.6190 ;
      RECT 0.8000 33.5080 55.6450 36.5090 ;
      RECT 0.8000 58.7120 55.6450 61.7130 ;
      RECT 0.0000 32.0330 55.6450 32.1080 ;
      RECT 0.8000 32.1220 54.8450 33.5080 ;
      RECT 0.0000 32.1080 54.8450 32.1220 ;
      RECT 0.8000 32.0070 54.8450 32.0190 ;
      RECT 0.8000 32.0190 55.6450 32.0330 ;
      RECT 0.0000 55.5690 1.5010 57.3590 ;
      RECT 0.8000 32.0190 54.8450 32.0330 ;
      RECT 0.0000 0.0000 20.5070 9.1790 ;
      RECT 0.0000 0.0000 20.5070 0.8000 ;
      RECT 0.8000 39.4630 54.8450 40.8490 ;
      RECT 0.8000 32.0330 54.8450 32.1080 ;
      RECT 0.8000 25.3280 54.8450 26.7140 ;
      RECT 0.8000 9.1800 54.8450 10.5790 ;
      RECT 0.0000 24.5380 54.8450 25.3280 ;
      RECT 0.0000 18.0990 54.8450 25.3280 ;
      RECT 0.0000 18.0990 54.8450 25.3280 ;
      RECT 0.0000 18.0990 54.8450 25.3280 ;
      RECT 0.0000 18.0990 55.6450 24.5380 ;
      RECT 0.0000 18.0460 54.8450 24.5380 ;
      RECT 0.0000 18.0460 54.8450 24.5380 ;
      RECT 0.0000 18.0460 54.8450 24.5380 ;
      RECT 0.0000 18.0460 54.8450 18.0990 ;
      RECT 0.0000 10.5800 55.6450 16.1860 ;
      RECT 0.8000 10.5800 54.8450 24.5380 ;
      RECT 0.8000 10.5800 54.8450 24.5380 ;
      RECT 0.8000 10.5800 54.8450 24.5380 ;
      RECT 0.8000 16.1920 54.8450 18.0460 ;
      RECT 0.8000 16.1860 55.6450 16.1920 ;
      RECT 0.8000 10.5800 55.6450 16.1920 ;
      RECT 0.8000 10.5800 55.6450 16.1920 ;
      RECT 0.8000 10.5800 55.6450 16.1920 ;
      RECT 0.8000 10.5790 55.6450 16.1860 ;
      RECT 0.8000 10.5790 55.6450 16.1860 ;
      RECT 0.8000 10.5790 55.6450 16.1860 ;
      RECT 0.8000 10.5790 55.6450 10.5800 ;
      RECT 0.0000 9.1790 54.8450 9.1800 ;
      RECT 0.0000 0.8000 54.8450 9.1800 ;
    LAYER PO ;
      RECT 0.0000 0.0000 55.6450 64.8190 ;
    LAYER M3 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 0.0000 53.7290 3.0010 54.0690 ;
      RECT 0.0000 55.6690 1.5010 57.2590 ;
      RECT 52.6440 58.8120 55.6450 58.8590 ;
      RECT 54.1440 55.6830 55.6450 57.2120 ;
      RECT 0.0000 18.1990 55.6450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 18.1990 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.0000 24.4380 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.0000 0.0000 20.4070 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 0.0000 26.8280 55.6450 29.8900 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 30.5190 54.7450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 30.5190 54.7450 33.6080 ;
      RECT 0.9000 26.8280 54.7450 33.6080 ;
      RECT 0.9000 29.8900 55.6450 30.5190 ;
      RECT 0.9000 26.8280 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
      RECT 0.0000 40.9630 55.6450 53.7290 ;
      RECT 0.9000 40.9630 54.7450 57.2120 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 40.9630 ;
      RECT 0.0000 58.8590 55.6450 64.8190 ;
      RECT 0.9000 55.6830 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
    LAYER M2 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 54.1440 55.6830 55.6450 57.2120 ;
      RECT 0.0000 55.6690 1.5010 57.2590 ;
      RECT 0.0000 53.7290 3.0010 54.0690 ;
      RECT 52.6440 58.8120 55.6450 58.8590 ;
      RECT 0.0000 18.1990 55.6450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 18.1990 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.0000 24.4380 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.0000 0.0000 20.4070 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 0.0000 26.8280 55.6450 29.8900 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 30.5190 54.7450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 30.5190 54.7450 33.6080 ;
      RECT 0.9000 26.8280 54.7450 33.6080 ;
      RECT 0.9000 29.8900 55.6450 30.5190 ;
      RECT 0.9000 26.8280 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
      RECT 0.0000 40.9630 55.6450 53.7290 ;
      RECT 0.9000 40.9630 54.7450 57.2120 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 40.9630 ;
      RECT 0.0000 58.8590 55.6450 64.8190 ;
      RECT 0.9000 55.6830 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
    LAYER M4 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.9000 30.5190 54.7450 33.6080 ;
      RECT 0.9000 26.8280 54.7450 33.6080 ;
      RECT 0.9000 29.8900 55.6450 30.5190 ;
      RECT 0.9000 26.8280 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 25.2280 54.7450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
      RECT 0.0000 40.9630 55.6450 53.7290 ;
      RECT 0.9000 40.9630 54.7450 57.2120 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 39.3630 54.7450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 40.9630 ;
      RECT 0.0000 58.8590 55.6450 64.8190 ;
      RECT 0.9000 55.6830 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 0.9000 54.0690 54.7450 64.8190 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 0.0000 53.7290 3.0010 54.0690 ;
      RECT 0.0000 55.6690 1.5010 57.2590 ;
      RECT 52.6440 58.8120 55.6450 58.8590 ;
      RECT 54.1440 55.6830 55.6450 57.2120 ;
      RECT 0.0000 18.1990 55.6450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 18.1990 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.0000 24.4380 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.0000 0.0000 20.4070 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 0.0000 26.8280 55.6450 29.8900 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 30.5190 54.7450 39.3490 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 55.6450 64.8190 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 55.6450 64.8190 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 55.6450 64.8190 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 55.6450 64.8190 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 55.6450 64.8190 ;
    LAYER M5 ;
      RECT 0.0000 63.8190 0.3650 64.8190 ;
      RECT 22.0070 0.0000 22.6950 0.9000 ;
      RECT 55.1650 63.8190 55.6450 64.8190 ;
      RECT 0.0000 55.6690 1.5010 57.2590 ;
      RECT 0.0000 51.0680 54.7450 54.0690 ;
      RECT 0.9000 58.8120 55.6450 61.8130 ;
      RECT 54.1440 55.6830 55.6450 57.2120 ;
      RECT 0.0000 39.3490 54.7450 39.3630 ;
      RECT 0.9000 39.3630 54.7450 40.9490 ;
      RECT 0.0000 0.0000 20.4070 9.0790 ;
      RECT 0.0000 0.0000 20.4070 0.9000 ;
      RECT 0.9000 9.0800 54.7450 10.6790 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 54.7450 39.3630 ;
      RECT 0.0000 33.6220 55.6450 39.3490 ;
      RECT 0.9000 33.6220 54.7450 40.9490 ;
      RECT 0.9000 33.6220 54.7450 40.9490 ;
      RECT 0.9000 33.6220 54.7450 40.9490 ;
      RECT 0.9000 33.6080 55.6450 39.3490 ;
      RECT 0.9000 33.6080 55.6450 33.6220 ;
      RECT 0.0000 10.6800 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 16.0860 ;
      RECT 0.9000 10.6790 55.6450 10.6800 ;
      RECT 0.9000 30.5190 54.7450 39.3490 ;
      RECT 0.9000 30.5190 54.7450 33.6080 ;
      RECT 0.0000 24.4380 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 54.7450 25.2280 ;
      RECT 0.0000 18.1990 55.6450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 24.4380 ;
      RECT 0.0000 18.1460 54.7450 18.1990 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 24.4380 ;
      RECT 0.9000 16.0920 54.7450 18.1460 ;
      RECT 0.9000 16.0860 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 10.6800 55.6450 16.0920 ;
      RECT 0.9000 29.8900 55.6450 30.5190 ;
      RECT 0.0000 26.8280 55.6450 29.8900 ;
      RECT 0.9000 26.8280 54.7450 33.6080 ;
      RECT 0.9000 26.8280 55.6450 30.5190 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 29.8900 ;
      RECT 0.9000 26.8140 55.6450 26.8280 ;
      RECT 0.9000 25.2280 54.7450 26.8140 ;
      RECT 0.9000 18.1990 54.7450 26.8140 ;
      RECT 0.9000 18.1990 54.7450 26.8140 ;
      RECT 0.9000 18.1990 54.7450 26.8140 ;
      RECT 0.0000 9.0790 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 54.7450 9.0800 ;
      RECT 0.0000 0.9000 55.6450 9.0790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 0.9000 0.9000 54.7450 10.6790 ;
      RECT 35.4390 0.0000 55.6450 9.0790 ;
      RECT 35.4390 0.0000 55.6450 0.9000 ;
      RECT 0.9000 55.6830 54.7450 57.2120 ;
      RECT 0.0000 58.8590 55.6450 63.8190 ;
      RECT 0.9000 55.6830 54.7450 58.8120 ;
      RECT 0.9000 57.2120 54.7450 57.2590 ;
      RECT 0.0000 40.9630 55.6450 53.7290 ;
      RECT 0.9000 55.6690 54.7450 58.8120 ;
      RECT 0.9000 55.6690 54.7450 58.8120 ;
      RECT 0.9000 55.6690 54.7450 58.8120 ;
      RECT 0.9000 55.6690 54.7450 58.8120 ;
      RECT 0.9000 55.6690 54.7450 58.8120 ;
      RECT 0.9000 54.0690 54.7450 58.8120 ;
      RECT 0.9000 54.0690 54.7450 58.8120 ;
      RECT 0.9000 54.0690 54.7450 58.8120 ;
      RECT 0.9000 54.0690 54.7450 58.8120 ;
      RECT 0.9000 54.0690 54.7450 58.8120 ;
      RECT 0.9000 55.6690 54.7450 55.6830 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 53.7290 ;
      RECT 0.9000 40.9490 55.6450 40.9630 ;
  END
END SRAMLP2RW32x4

MACRO SRAMLP2RW32x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 69.453 BY 67.414 ;
  SYMMETRY X Y R90 ;

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.9050 0.0000 32.1050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.9050 0.0000 32.1050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.9050 0.0000 32.1050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.9050 0.0000 32.1050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[2]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.5800 0.0000 42.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.5800 0.0000 42.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.5800 0.0000 42.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.5800 0.0000 42.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.5800 0.0000 42.7800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[2]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2120 0.0000 41.4120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2120 0.0000 41.4120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2120 0.0000 41.4120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2120 0.0000 41.4120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2120 0.0000 41.4120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[4]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.6190 0.0000 44.8190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.6190 0.0000 44.8190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.6190 0.0000 44.8190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.6190 0.0000 44.8190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.6190 0.0000 44.8190 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.2510 0.0000 43.4510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.2510 0.0000 43.4510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.2510 0.0000 43.4510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.2510 0.0000 43.4510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.2510 0.0000 43.4510 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[2]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3160 0.0000 45.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3160 0.0000 45.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3160 0.0000 45.5160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3160 0.0000 45.5160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3160 0.0000 45.5160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[5]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.9480 0.0000 44.1480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.9480 0.0000 44.1480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.9480 0.0000 44.1480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.9480 0.0000 44.1480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.9480 0.0000 44.1480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[3]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.9870 0.0000 46.1870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.9870 0.0000 46.1870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.9870 0.0000 46.1870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.9870 0.0000 46.1870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.9870 0.0000 46.1870 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[5]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 9.8550 69.4530 10.0550 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 9.8550 69.4530 10.0550 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 9.8550 69.4530 10.0550 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 9.8550 69.4530 10.0550 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 9.8550 69.4530 10.0550 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8550 0.2000 10.0550 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8550 0.2000 10.0550 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8550 0.2000 10.0550 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8550 0.2000 10.0550 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8550 0.2000 10.0550 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 60.4620 69.4530 60.6620 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 60.4620 69.4530 60.6620 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 60.4620 69.4530 60.6620 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 60.4620 69.4530 60.6620 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 60.4620 69.4530 60.6620 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 57.2360 0.2000 57.4360 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 57.2360 0.2000 57.4360 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 57.2360 0.2000 57.4360 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 57.2360 0.2000 57.4360 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 57.2360 0.2000 57.4360 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 60.4220 0.2000 60.6220 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 60.4220 0.2000 60.6220 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 60.4220 0.2000 60.6220 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 60.4220 0.2000 60.6220 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 60.4220 0.2000 60.6220 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.1050 0.0000 22.3050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.1050 0.0000 22.3050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.1050 0.0000 22.3050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.1050 0.0000 22.3050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.1050 0.0000 22.3050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.4810 0.0000 46.6810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.4810 0.0000 46.6810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.4810 0.0000 46.6810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.4810 0.0000 46.6810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.4810 0.0000 46.6810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 28.2140 69.4530 28.4140 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 28.2140 69.4530 28.4140 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 28.2140 69.4530 28.4140 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 28.2140 69.4530 28.4140 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 28.2140 69.4530 28.4140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.2140 0.2000 28.4140 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 28.2140 0.2000 28.4140 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 28.2140 0.2000 28.4140 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 28.2140 0.2000 28.4140 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 28.2140 0.2000 28.4140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[4]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.1690 0.0000 29.3690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.1690 0.0000 29.3690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.1690 0.0000 29.3690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.1690 0.0000 29.3690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.1690 0.0000 29.3690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[6]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.5370 0.0000 30.7370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.5370 0.0000 30.7370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.5370 0.0000 30.7370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.5370 0.0000 30.7370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.5370 0.0000 30.7370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[4]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.8660 0.0000 30.0660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.8660 0.0000 30.0660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.8660 0.0000 30.0660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.8660 0.0000 30.0660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.8660 0.0000 30.0660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[4]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.2340 0.0000 31.4340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.2340 0.0000 31.4340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.2340 0.0000 31.4340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.2340 0.0000 31.4340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.2340 0.0000 31.4340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[2]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.2730 0.0000 33.4730 0.2000 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.9050 0.0000 32.1050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.2730 0.0000 33.4730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.2730 0.0000 33.4730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.2730 0.0000 33.4730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.2730 0.0000 33.4730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[3]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.6020 0.0000 32.8020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.6020 0.0000 32.8020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.6020 0.0000 32.8020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.6020 0.0000 32.8020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.6020 0.0000 32.8020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[3]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.6410 0.0000 34.8410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.6410 0.0000 34.8410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.6410 0.0000 34.8410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.6410 0.0000 34.8410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.6410 0.0000 34.8410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[5]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.9700 0.0000 34.1700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.9700 0.0000 34.1700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.9700 0.0000 34.1700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.9700 0.0000 34.1700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.9700 0.0000 34.1700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[5]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4110 0.0000 36.6110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4110 0.0000 36.6110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4110 0.0000 36.6110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4110 0.0000 36.6110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4110 0.0000 36.6110 0.2000 ;
    END
    ANTENNADIFFAREA 1.9074 LAYER M3 ;
    ANTENNADIFFAREA 1.9074 LAYER M4 ;
    ANTENNADIFFAREA 1.9074 LAYER M5 ;
    ANTENNADIFFAREA 1.9074 LAYER M6 ;
    ANTENNADIFFAREA 1.9074 LAYER M7 ;
    ANTENNADIFFAREA 1.9074 LAYER M8 ;
    ANTENNADIFFAREA 1.9074 LAYER M9 ;
    ANTENNADIFFAREA 1.9074 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.2844 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.09504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.09504 LAYER M3 ;
    ANTENNAMAXAREACAR 22.04699 LAYER M3 ;
    ANTENNAGATEAREA 0.2844 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M4 ;
    ANTENNAMAXAREACAR 26.31122 LAYER M4 ;
    ANTENNAGATEAREA 0.2844 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M5 ;
    ANTENNAMAXAREACAR 30.57542 LAYER M5 ;
    ANTENNAGATEAREA 0.2844 LAYER M6 ;
    ANTENNAGATEAREA 0.2844 LAYER M7 ;
    ANTENNAGATEAREA 0.2844 LAYER M8 ;
    ANTENNAGATEAREA 0.2844 LAYER M9 ;
    ANTENNAGATEAREA 0.2844 LAYER MRDL ;
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.7400 0.0000 35.9400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.7400 0.0000 35.9400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.7400 0.0000 35.9400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.7400 0.0000 35.9400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.7400 0.0000 35.9400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[0]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1080 0.0000 37.3080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1080 0.0000 37.3080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1080 0.0000 37.3080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1080 0.0000 37.3080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1080 0.0000 37.3080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[7]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.1470 0.0000 39.3470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.1470 0.0000 39.3470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.1470 0.0000 39.3470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.1470 0.0000 39.3470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.1470 0.0000 39.3470 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[1]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.7790 0.0000 37.9790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.7790 0.0000 37.9790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.7790 0.0000 37.9790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.7790 0.0000 37.9790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.7790 0.0000 37.9790 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[7]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8440 0.0000 40.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.8440 0.0000 40.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.8440 0.0000 40.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.8440 0.0000 40.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.8440 0.0000 40.0440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[6]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.4760 0.0000 38.6760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.4760 0.0000 38.6760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.4760 0.0000 38.6760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.4760 0.0000 38.6760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.4760 0.0000 38.6760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[1]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.8830 0.0000 42.0830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.8830 0.0000 42.0830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.8830 0.0000 42.0830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.8830 0.0000 42.0830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.8830 0.0000 42.0830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[4]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5150 0.0000 40.7150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5150 0.0000 40.7150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5150 0.0000 40.7150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5150 0.0000 40.7150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5150 0.0000 40.7150 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[6]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 38.1190 69.4530 38.3190 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 38.1190 69.4530 38.3190 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 38.1190 69.4530 38.3190 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 38.1190 69.4530 38.3190 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 38.1190 69.4530 38.3190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 45.4190 69.4530 45.6190 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 45.4190 69.4530 45.6190 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 45.4190 69.4530 45.6190 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 45.4190 69.4530 45.6190 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 45.4190 69.4530 45.6190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 46.9410 69.4530 47.1410 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 46.9410 69.4530 47.1410 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 46.9410 69.4530 47.1410 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 46.9410 69.4530 47.1410 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 46.9410 69.4530 47.1410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 54.2340 69.4530 54.4340 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 54.2340 69.4530 54.4340 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 54.2340 69.4530 54.4340 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 54.2340 69.4530 54.4340 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 54.2340 69.4530 54.4340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 56.9080 69.4530 57.1080 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 56.9080 69.4530 57.1080 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 56.9080 69.4530 57.1080 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 56.9080 69.4530 57.1080 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 56.9080 69.4530 57.1080 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8670 0.2000 17.0670 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8670 0.2000 17.0670 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8670 0.2000 17.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8670 0.2000 17.0670 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8670 0.2000 17.0670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4020 0.2000 17.6020 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4020 0.2000 17.6020 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4020 0.2000 17.6020 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4020 0.2000 17.6020 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4020 0.2000 17.6020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE2

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 38.1190 0.2000 38.3190 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 38.1190 0.2000 38.3190 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 38.1190 0.2000 38.3190 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 38.1190 0.2000 38.3190 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 38.1190 0.2000 38.3190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.4190 0.2000 45.6190 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 45.4190 0.2000 45.6190 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 45.4190 0.2000 45.6190 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 45.4190 0.2000 45.6190 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 45.4190 0.2000 45.6190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 46.9400 0.2000 47.1400 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 46.9400 0.2000 47.1400 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 46.9400 0.2000 47.1400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 46.9400 0.2000 47.1400 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 46.9400 0.2000 47.1400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 54.2340 0.2000 54.4340 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 54.2340 0.2000 54.4340 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 54.2340 0.2000 54.4340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 54.2340 0.2000 54.4340 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 54.2340 0.2000 54.4340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.4330 0.0000 26.6330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.4330 0.0000 26.6330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.4330 0.0000 26.6330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.4330 0.0000 26.6330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.4330 0.0000 26.6330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[7]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.0650 0.0000 25.2650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.0650 0.0000 25.2650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.0650 0.0000 25.2650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.0650 0.0000 25.2650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.0650 0.0000 25.2650 0.2000 ;
    END
    ANTENNADIFFAREA 1.84416 LAYER M3 ;
    ANTENNADIFFAREA 1.84416 LAYER M4 ;
    ANTENNADIFFAREA 1.84416 LAYER M5 ;
    ANTENNADIFFAREA 1.84416 LAYER M6 ;
    ANTENNADIFFAREA 1.84416 LAYER M7 ;
    ANTENNADIFFAREA 1.84416 LAYER M8 ;
    ANTENNADIFFAREA 1.84416 LAYER M9 ;
    ANTENNADIFFAREA 1.84416 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.1716 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.09504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.09504 LAYER M3 ;
    ANTENNAMAXAREACAR 24.99795 LAYER M3 ;
    ANTENNAGATEAREA 0.1716 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M4 ;
    ANTENNAMAXAREACAR 32.06535 LAYER M4 ;
    ANTENNAGATEAREA 0.1716 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1.2128 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2128 LAYER M5 ;
    ANTENNAMAXAREACAR 39.13268 LAYER M5 ;
    ANTENNAGATEAREA 0.1716 LAYER M6 ;
    ANTENNAGATEAREA 0.1716 LAYER M7 ;
    ANTENNAGATEAREA 0.1716 LAYER M8 ;
    ANTENNAGATEAREA 0.1716 LAYER M9 ;
    ANTENNAGATEAREA 0.1716 LAYER MRDL ;
  END O2[0]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.3940 0.0000 24.5940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.3940 0.0000 24.5940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.3940 0.0000 24.5940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.3940 0.0000 24.5940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.3940 0.0000 24.5940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[0]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.7620 0.0000 25.9620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.7620 0.0000 25.9620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.7620 0.0000 25.9620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.7620 0.0000 25.9620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.7620 0.0000 25.9620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[7]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.8010 0.0000 28.0010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.8010 0.0000 28.0010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.8010 0.0000 28.0010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.8010 0.0000 28.0010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.8010 0.0000 28.0010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[1]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.1300 0.0000 27.3300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.1300 0.0000 27.3300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.1300 0.0000 27.3300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.1300 0.0000 27.3300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.1300 0.0000 27.3300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[1]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.4980 0.0000 28.6980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.4980 0.0000 28.6980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.4980 0.0000 28.6980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.4980 0.0000 28.6980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.4980 0.0000 28.6980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[6]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 16.8660 69.4530 17.0660 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 16.8660 69.4530 17.0660 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 16.8660 69.4530 17.0660 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 16.8660 69.4530 17.0660 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 16.8660 69.4530 17.0660 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.53692 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.53692 LAYER M4 ;
    ANTENNAMAXAREACAR 17.81934 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 21.96024 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 17.3260 69.4530 17.5260 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 17.3260 69.4530 17.5260 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 17.3260 69.4530 17.5260 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 17.3260 69.4530 17.5260 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 17.3260 69.4530 17.5260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15634 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.1128 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.85044 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85044 LAYER M4 ;
    ANTENNAMAXAREACAR 24.24627 LAYER M4 ;
    ANTENNAGATEAREA 0.1128 LAYER M5 ;
    ANTENNAGATEAREA 0.1128 LAYER M6 ;
    ANTENNAGATEAREA 0.1128 LAYER M7 ;
    ANTENNAGATEAREA 0.1128 LAYER M8 ;
    ANTENNAGATEAREA 0.1128 LAYER M9 ;
    ANTENNAGATEAREA 0.1128 LAYER MRDL ;
  END CE1

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.2530 57.2480 69.4530 57.4480 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.2530 57.2480 69.4530 57.4480 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.2530 57.2480 69.4530 57.4480 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.2530 57.2480 69.4530 57.4480 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.2530 57.2480 69.4530 57.4480 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
  END DS1

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 61.0370 67.1140 61.3370 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.1370 67.1140 60.4360 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.7370 67.1140 19.0360 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.6370 67.1140 19.9370 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.8360 67.1140 9.1370 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.9360 67.1140 8.2370 67.4140 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 119.6073 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 119.6073 LAYER M5 ;
  END VDDL

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 61.9360 67.1140 62.2350 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.8360 67.1140 63.1350 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.9370 67.1140 17.2370 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.0360 67.1140 16.3360 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.2360 67.1140 5.5360 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.1370 67.1140 6.4360 67.4140 ;
    END
    ANTENNADIFFAREA 11.07611 LAYER M5 ;
    ANTENNADIFFAREA 11.07611 LAYER M6 ;
    ANTENNADIFFAREA 11.07611 LAYER M7 ;
    ANTENNADIFFAREA 11.07611 LAYER M8 ;
    ANTENNADIFFAREA 11.07611 LAYER M9 ;
    ANTENNADIFFAREA 11.07611 LAYER MRDL ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 119.6076 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 119.6076 LAYER M5 ;
    ANTENNAMAXAREACAR 2784.928 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 7.4870 67.1140 7.7870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.4870 67.1140 16.7860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.2860 67.1140 18.5870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.1860 67.1140 19.4870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.0860 67.1140 20.3870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.3870 67.1140 8.6860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.9870 67.1140 12.2870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.7860 67.1140 14.0860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.8870 67.1140 13.1860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.6870 67.1140 14.9870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.5860 67.1140 15.8860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.3860 67.1140 17.6860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.6860 67.1140 23.9870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.3860 67.1140 26.6870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.8870 67.1140 22.1870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.7860 67.1140 23.0860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.9870 67.1140 21.2870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.2860 67.1140 27.5860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.4870 67.1140 25.7860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.5870 67.1140 24.8870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.6860 67.1140 32.9870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.5860 67.1140 33.8870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.1870 67.1140 28.4870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.7870 67.1140 32.0860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.8870 67.1140 31.1860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.9870 67.1140 30.2870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.0860 67.1140 29.3860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.3870 67.1140 35.6860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.4870 67.1140 34.7870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.1860 67.1140 37.4870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.0860 67.1140 38.3870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.5870 67.1140 42.8880 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.2870 67.1140 36.5860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.9860 67.1140 39.2860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.8860 67.1140 40.1860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.7870 67.1140 41.0870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.6860 67.1140 41.9850 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.0870 67.1140 47.3880 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.4860 67.1140 43.7860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.3860 67.1140 44.6860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.2870 67.1140 45.5870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.1860 67.1140 46.4850 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.9860 67.1140 48.2860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.7870 67.1140 50.0870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.8860 67.1140 49.1860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.5870 67.1140 51.8880 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.6860 67.1140 50.9850 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.8850 67.1140 67.1850 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.0860 67.1140 65.3860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.4870 67.1140 61.7870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.8870 67.1140 58.1870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.2870 67.1140 54.5870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.4860 67.1140 52.7860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.9850 67.1140 66.2850 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.1850 67.1140 64.4850 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.2860 67.1140 63.5860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.3860 67.1140 62.6860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.5860 67.1140 60.8860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.6860 67.1140 59.9860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.7860 67.1140 59.0860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.9860 67.1140 57.2860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.0860 67.1140 56.3860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.1860 67.1140 55.4860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.3860 67.1140 53.6860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.0840 67.1140 2.3840 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.5860 67.1140 6.8870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.6860 67.1140 5.9870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.0860 67.1140 11.3870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.1860 67.1140 10.4870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.8870 67.1140 4.1870 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.9860 67.1140 3.2860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.7860 67.1140 5.0860 67.4140 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.2870 67.1140 9.5860 67.4140 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 53.6340 68.6530 61.2220 ;
      RECT 0.8000 53.6340 68.6530 61.2220 ;
      RECT 0.8000 59.8220 68.6530 59.8620 ;
      RECT 0.8000 58.0480 68.6530 59.8220 ;
      RECT 0.8000 56.6360 68.6530 59.8220 ;
      RECT 0.8000 56.6360 68.6530 59.8220 ;
      RECT 0.8000 56.6360 68.6530 59.8220 ;
      RECT 0.8000 56.3080 68.6530 59.8220 ;
      RECT 0.8000 56.3080 68.6530 59.8220 ;
      RECT 0.8000 56.3080 68.6530 59.8220 ;
      RECT 0.8000 58.0360 68.6530 58.0480 ;
      RECT 0.8000 56.6360 68.6530 58.0360 ;
      RECT 0.8000 56.3080 68.6530 56.6360 ;
      RECT 0.8000 53.6340 68.6530 56.6360 ;
      RECT 0.8000 53.6340 68.6530 56.6360 ;
      RECT 0.8000 55.0340 68.6530 56.3080 ;
      RECT 0.0000 10.6550 69.4530 16.2660 ;
      RECT 0.8000 9.2550 68.6530 10.6550 ;
      RECT 0.8000 0.8000 68.6530 10.6550 ;
      RECT 0.0000 18.2020 69.4530 27.6140 ;
      RECT 0.0000 16.2660 68.6530 16.2670 ;
      RECT 0.0000 10.6550 68.6530 16.2670 ;
      RECT 0.0000 10.6550 68.6530 16.2670 ;
      RECT 0.0000 10.6550 68.6530 16.2670 ;
      RECT 0.8000 27.6140 68.6530 29.0140 ;
      RECT 0.8000 18.2020 68.6530 29.0140 ;
      RECT 0.8000 18.1260 69.4530 27.6140 ;
      RECT 0.8000 18.1260 69.4530 27.6140 ;
      RECT 0.8000 18.1260 69.4530 27.6140 ;
      RECT 0.8000 16.2670 68.6530 27.6140 ;
      RECT 0.8000 16.2670 68.6530 27.6140 ;
      RECT 0.8000 16.2670 68.6530 27.6140 ;
      RECT 0.8000 18.1260 69.4530 18.2020 ;
      RECT 0.8000 16.2670 68.6530 18.1260 ;
      RECT 0.0000 46.2190 0.8000 46.3400 ;
      RECT 68.6530 55.0340 69.4530 56.3080 ;
      RECT 22.9050 0.0000 23.7940 0.8000 ;
      RECT 0.0000 55.0340 1.5010 56.6360 ;
      RECT 0.0000 58.0360 1.5010 59.8220 ;
      RECT 67.9520 58.0480 69.4530 59.8620 ;
      RECT 68.6530 46.2190 69.4530 46.3410 ;
      RECT 0.8000 46.3410 68.6530 47.7400 ;
      RECT 0.8000 46.3400 68.6530 46.3410 ;
      RECT 0.8000 46.2190 68.6530 46.3400 ;
      RECT 0.8000 44.8190 68.6530 46.2190 ;
      RECT 0.0000 0.0000 21.5050 9.2550 ;
      RECT 0.0000 0.8000 69.4530 9.2550 ;
      RECT 0.0000 0.0000 21.5050 0.8000 ;
      RECT 47.2810 0.0000 69.4530 9.2550 ;
      RECT 47.2810 0.0000 69.4530 0.8000 ;
      RECT 0.0000 38.9190 69.4530 44.8190 ;
      RECT 0.0000 29.0140 69.4530 37.5190 ;
      RECT 0.8000 37.5190 68.6530 38.9190 ;
      RECT 0.8000 29.0140 68.6530 38.9190 ;
      RECT 0.0000 61.2620 69.4530 67.4140 ;
      RECT 0.0000 61.2220 68.6530 67.4140 ;
      RECT 0.0000 61.2220 68.6530 67.4140 ;
      RECT 0.0000 61.2220 68.6530 67.4140 ;
      RECT 0.0000 61.2220 68.6530 67.4140 ;
      RECT 0.0000 61.2220 68.6530 61.2620 ;
      RECT 0.8000 59.8620 68.6530 61.2220 ;
      RECT 0.0000 47.7410 69.4530 53.6340 ;
      RECT 0.0000 47.7400 68.6530 47.7410 ;
      RECT 0.8000 53.6340 68.6530 55.0340 ;
      RECT 0.8000 47.7410 68.6530 55.0340 ;
      RECT 0.8000 47.7410 68.6530 55.0340 ;
      RECT 0.8000 47.7410 68.6530 55.0340 ;
      RECT 0.8000 47.7410 68.6530 55.0340 ;
      RECT 0.8000 58.0480 68.6530 67.4140 ;
      RECT 0.8000 58.0480 68.6530 67.4140 ;
      RECT 0.8000 58.0480 68.6530 61.2220 ;
      RECT 0.8000 58.0480 68.6530 61.2220 ;
      RECT 0.8000 58.0480 68.6530 61.2220 ;
      RECT 0.8000 58.0480 68.6530 61.2220 ;
      RECT 0.8000 58.0480 68.6530 61.2220 ;
      RECT 0.8000 58.0480 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
      RECT 0.8000 56.6360 68.6530 61.2220 ;
    LAYER PO ;
      RECT 0.0000 0.0000 69.4530 67.4140 ;
    LAYER M3 ;
      RECT 0.9000 58.1360 68.5530 58.1480 ;
      RECT 0.9000 56.5360 68.5530 58.1360 ;
      RECT 0.9000 56.2080 68.5530 56.5360 ;
      RECT 0.9000 55.1340 68.5530 56.2080 ;
      RECT 0.9000 53.5340 68.5530 55.1340 ;
      RECT 0.9000 44.7190 68.5530 47.8400 ;
      RECT 0.9000 37.4190 68.5530 39.0190 ;
      RECT 0.9000 27.5140 68.5530 29.1140 ;
      RECT 0.9000 18.2260 69.4530 27.5140 ;
      RECT 0.9000 18.2260 69.4530 18.3020 ;
      RECT 0.9000 16.1670 68.5530 18.2260 ;
      RECT 0.9000 9.1550 68.5530 10.7550 ;
      RECT 47.3810 0.0000 69.4530 9.1550 ;
      RECT 47.3810 0.0000 69.4530 0.9000 ;
      RECT 0.0000 61.3620 69.4530 67.4140 ;
      RECT 0.0000 61.3220 68.5530 67.4140 ;
      RECT 0.0000 61.3220 68.5530 61.3620 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 59.7620 68.5530 61.3220 ;
      RECT 23.0050 0.0000 23.6940 0.9000 ;
      RECT 0.0000 58.1360 1.5010 59.7220 ;
      RECT 0.0000 55.1340 0.9000 56.5360 ;
      RECT 67.9520 58.1480 69.4530 59.7620 ;
      RECT 68.5530 55.1340 69.4530 56.2080 ;
      RECT 0.0000 47.8410 69.4530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 47.8410 ;
      RECT 0.0000 39.0190 69.4530 44.7190 ;
      RECT 0.0000 29.1140 69.4530 37.4190 ;
      RECT 0.0000 18.3020 69.4530 27.5140 ;
      RECT 0.0000 16.1660 68.5530 16.1670 ;
      RECT 0.0000 10.7550 68.5530 16.1670 ;
      RECT 0.0000 10.7550 69.4530 16.1660 ;
      RECT 0.0000 0.0000 21.4050 9.1550 ;
      RECT 0.0000 0.9000 69.4530 9.1550 ;
      RECT 0.0000 0.0000 21.4050 0.9000 ;
      RECT 0.9000 59.7220 68.5530 59.7620 ;
      RECT 0.9000 58.1480 68.5530 59.7220 ;
    LAYER M2 ;
      RECT 0.0000 55.1340 0.9000 56.5360 ;
      RECT 68.5530 55.1340 69.4530 56.2080 ;
      RECT 23.0050 0.0000 23.6940 0.9000 ;
      RECT 0.0000 58.1360 1.5010 59.7220 ;
      RECT 67.9520 58.1480 69.4530 59.7620 ;
      RECT 0.0000 47.8410 69.4530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 47.8410 ;
      RECT 0.0000 39.0190 69.4530 44.7190 ;
      RECT 0.0000 29.1140 69.4530 37.4190 ;
      RECT 0.0000 18.3020 69.4530 27.5140 ;
      RECT 0.0000 16.1660 68.5530 16.1670 ;
      RECT 0.0000 10.7550 68.5530 16.1670 ;
      RECT 0.0000 10.7550 69.4530 16.1660 ;
      RECT 0.0000 0.0000 21.4050 9.1550 ;
      RECT 0.0000 0.9000 69.4530 9.1550 ;
      RECT 0.0000 0.0000 21.4050 0.9000 ;
      RECT 0.9000 59.7220 68.5530 59.7620 ;
      RECT 0.9000 58.1480 68.5530 59.7220 ;
      RECT 0.9000 58.1360 68.5530 58.1480 ;
      RECT 0.9000 56.5360 68.5530 58.1360 ;
      RECT 0.9000 56.2080 68.5530 56.5360 ;
      RECT 0.9000 55.1340 68.5530 56.2080 ;
      RECT 0.9000 53.5340 68.5530 55.1340 ;
      RECT 0.9000 44.7190 68.5530 47.8400 ;
      RECT 0.9000 37.4190 68.5530 39.0190 ;
      RECT 0.9000 27.5140 68.5530 29.1140 ;
      RECT 0.9000 18.2260 69.4530 27.5140 ;
      RECT 0.9000 18.2260 69.4530 18.3020 ;
      RECT 0.9000 16.1670 68.5530 18.2260 ;
      RECT 0.9000 9.1550 68.5530 10.7550 ;
      RECT 47.3810 0.0000 69.4530 9.1550 ;
      RECT 47.3810 0.0000 69.4530 0.9000 ;
      RECT 0.0000 61.3620 69.4530 67.4140 ;
      RECT 0.0000 61.3220 68.5530 67.4140 ;
      RECT 0.0000 61.3220 68.5530 61.3620 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 59.7620 68.5530 61.3220 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 69.4530 67.4140 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 69.4530 67.4140 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 69.4530 67.4140 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 69.4530 67.4140 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 69.4530 67.4140 ;
    LAYER M5 ;
      RECT 0.0000 66.4140 1.3840 67.4140 ;
      RECT 23.0050 0.0000 23.6940 0.9000 ;
      RECT 67.8850 66.4140 69.4530 67.4140 ;
      RECT 0.0000 58.1360 1.5010 59.7220 ;
      RECT 0.0000 55.1340 0.9000 56.5360 ;
      RECT 67.8850 65.9130 69.4530 67.4140 ;
      RECT 67.9520 58.1480 69.4530 59.7620 ;
      RECT 68.5530 55.1340 69.4530 56.2080 ;
      RECT 0.0000 47.8410 69.4530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 47.8410 ;
      RECT 0.0000 39.0190 69.4530 44.7190 ;
      RECT 0.0000 29.1140 69.4530 37.4190 ;
      RECT 0.0000 18.3020 69.4530 27.5140 ;
      RECT 0.0000 16.1660 68.5530 16.1670 ;
      RECT 0.0000 10.7550 68.5530 16.1670 ;
      RECT 0.0000 10.7550 69.4530 16.1660 ;
      RECT 0.0000 0.0000 21.4050 9.1550 ;
      RECT 0.0000 0.9000 69.4530 9.1550 ;
      RECT 0.0000 0.0000 21.4050 0.9000 ;
      RECT 0.9000 59.7220 68.5530 59.7620 ;
      RECT 0.9000 58.1480 68.5530 59.7220 ;
      RECT 0.9000 58.1360 68.5530 58.1480 ;
      RECT 0.9000 56.5360 68.5530 58.1360 ;
      RECT 0.9000 56.2080 68.5530 56.5360 ;
      RECT 0.9000 55.1340 68.5530 56.2080 ;
      RECT 0.9000 53.5340 68.5530 55.1340 ;
      RECT 0.9000 44.7190 68.5530 47.8400 ;
      RECT 0.9000 37.4190 68.5530 39.0190 ;
      RECT 0.9000 27.5140 68.5530 29.1140 ;
      RECT 0.9000 18.2260 69.4530 27.5140 ;
      RECT 0.9000 18.2260 69.4530 18.3020 ;
      RECT 0.9000 16.1670 68.5530 18.2260 ;
      RECT 0.9000 9.1550 68.5530 10.7550 ;
      RECT 47.3810 0.0000 69.4530 9.1550 ;
      RECT 47.3810 0.0000 69.4530 0.9000 ;
      RECT 0.0000 61.3620 69.4530 66.4140 ;
      RECT 0.0000 61.3220 68.5530 66.4140 ;
      RECT 0.0000 61.3220 68.5530 61.3620 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 0.9000 68.5530 66.4140 ;
      RECT 0.9000 59.7620 68.5530 61.3220 ;
    LAYER M4 ;
      RECT 23.0050 0.0000 23.6940 0.9000 ;
      RECT 0.0000 58.1360 1.5010 59.7220 ;
      RECT 0.0000 55.1340 0.9000 56.5360 ;
      RECT 67.9520 58.1480 69.4530 59.7620 ;
      RECT 68.5530 55.1340 69.4530 56.2080 ;
      RECT 0.0000 47.8410 69.4530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 53.5340 ;
      RECT 0.0000 47.8400 68.5530 47.8410 ;
      RECT 0.0000 39.0190 69.4530 44.7190 ;
      RECT 0.0000 29.1140 69.4530 37.4190 ;
      RECT 0.0000 18.3020 69.4530 27.5140 ;
      RECT 0.0000 16.1660 68.5530 16.1670 ;
      RECT 0.0000 10.7550 68.5530 16.1670 ;
      RECT 0.0000 10.7550 69.4530 16.1660 ;
      RECT 0.0000 0.0000 21.4050 9.1550 ;
      RECT 0.0000 0.9000 69.4530 9.1550 ;
      RECT 0.0000 0.0000 21.4050 0.9000 ;
      RECT 0.9000 59.7220 68.5530 59.7620 ;
      RECT 0.9000 58.1480 68.5530 59.7220 ;
      RECT 0.9000 58.1360 68.5530 58.1480 ;
      RECT 0.9000 56.5360 68.5530 58.1360 ;
      RECT 0.9000 56.2080 68.5530 56.5360 ;
      RECT 0.9000 55.1340 68.5530 56.2080 ;
      RECT 0.9000 53.5340 68.5530 55.1340 ;
      RECT 0.9000 44.7190 68.5530 47.8400 ;
      RECT 0.9000 37.4190 68.5530 39.0190 ;
      RECT 0.9000 27.5140 68.5530 29.1140 ;
      RECT 0.9000 18.2260 69.4530 27.5140 ;
      RECT 0.9000 18.2260 69.4530 18.3020 ;
      RECT 0.9000 16.1670 68.5530 18.2260 ;
      RECT 0.9000 9.1550 68.5530 10.7550 ;
      RECT 47.3810 0.0000 69.4530 9.1550 ;
      RECT 47.3810 0.0000 69.4530 0.9000 ;
      RECT 0.0000 61.3620 69.4530 67.4140 ;
      RECT 0.0000 61.3220 68.5530 67.4140 ;
      RECT 0.0000 61.3220 68.5530 61.3620 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 0.9000 68.5530 67.4140 ;
      RECT 0.9000 59.7620 68.5530 61.3220 ;
  END
END SRAMLP2RW32x8

MACRO SRAMLP2RW32x16
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 93.479 BY 73.52 ;
  SYMMETRY X Y R90 ;

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.9000 0.0000 70.1000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.9000 0.0000 70.1000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.9000 0.0000 70.1000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.9000 0.0000 70.1000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.9000 0.0000 70.1000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 42.6960 0.2000 42.8960 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 50.0630 0.2000 50.2630 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 51.2600 0.2000 51.4600 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 58.4900 0.2000 58.6900 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 42.6960 0.2000 42.8960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 50.0630 0.2000 50.2630 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 51.2600 0.2000 51.4600 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 58.4900 0.2000 58.6900 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 42.6960 0.2000 42.8960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 50.0630 0.2000 50.2630 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 51.2600 0.2000 51.4600 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 58.4900 0.2000 58.6900 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 42.6960 0.2000 42.8960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 50.0630 0.2000 50.2630 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 51.2600 0.2000 51.4600 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 58.4900 0.2000 58.6900 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 58.4900 0.2000 58.6900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 58.4900 93.4790 58.6900 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 58.4900 93.4790 58.6900 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 58.4900 93.4790 58.6900 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 58.4900 93.4790 58.6900 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 58.4900 93.4790 58.6900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 17.2900 93.4790 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 17.2900 93.4790 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 17.2900 93.4790 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 17.2900 93.4790 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 17.2900 93.4790 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 16.8310 93.4790 17.0310 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 16.8310 93.4790 17.0310 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 16.8310 93.4790 17.0310 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 16.8310 93.4790 17.0310 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 16.8310 93.4790 17.0310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB1

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 32.4850 93.4790 32.6850 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 32.4850 93.4790 32.6850 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 32.4850 93.4790 32.6850 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 32.4850 93.4790 32.6850 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 32.4850 93.4790 32.6850 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 49.4650 93.4790 49.6650 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 49.4650 93.4790 49.6650 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 49.4650 93.4790 49.6650 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 49.4650 93.4790 49.6650 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 49.4650 93.4790 49.6650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 42.6130 93.4790 42.8130 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 42.6130 93.4790 42.8130 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 42.6130 93.4790 42.8130 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 42.6130 93.4790 42.8130 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 42.6130 93.4790 42.8130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 51.2600 93.4790 51.4600 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 51.2600 93.4790 51.4600 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 51.2600 93.4790 51.4600 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 51.2600 93.4790 51.4600 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 51.2600 93.4790 51.4600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 11.2640 73.2200 11.5640 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1650 73.2200 12.4650 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.3640 73.2200 91.6640 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3630 73.2200 1.6630 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.2660 73.2200 92.5650 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2620 73.2200 2.5620 73.5200 ;
    END
    ANTENNADIFFAREA 10.95167 LAYER M5 ;
    ANTENNADIFFAREA 10.95167 LAYER M6 ;
    ANTENNADIFFAREA 10.95167 LAYER M7 ;
    ANTENNADIFFAREA 10.95167 LAYER M8 ;
    ANTENNADIFFAREA 10.95167 LAYER M9 ;
    ANTENNADIFFAREA 10.95167 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 130.6575 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 130.6575 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 5.4140 73.2200 5.7140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.5140 73.2200 4.8140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6140 73.2200 3.9140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7140 73.2200 3.0140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.8140 73.2200 2.1140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.9150 73.2200 10.2150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.0140 73.2200 9.3140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.1150 73.2200 8.4150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.2140 73.2200 7.5140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.3150 73.2200 6.6150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.4150 73.2200 14.7150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.5140 73.2200 13.8140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6140 73.2200 12.9140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7150 73.2200 12.0150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.8150 73.2200 11.1150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.8150 73.2200 20.1150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.9150 73.2200 19.2150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0140 73.2200 18.3140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1150 73.2200 17.4150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.2150 73.2200 16.5150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.3150 73.2200 15.6150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.5150 73.2200 22.8150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.4160 73.2200 23.7160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.7160 73.2200 21.0160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.3150 73.2200 24.6140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.6150 73.2200 21.9150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.9150 73.2200 28.2150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.8160 73.2200 29.1160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.1150 73.2200 26.4150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.2160 73.2200 25.5170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.0150 73.2200 27.3150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.2150 73.2200 34.5140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.4150 73.2200 32.7150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.7150 73.2200 30.0140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.5150 73.2200 31.8150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.3150 73.2200 33.6150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.6160 73.2200 30.9170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.7150 73.2200 39.0150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.9150 73.2200 37.2150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.8160 73.2200 38.1160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.0150 73.2200 36.3150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.1160 73.2200 35.4170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.5160 73.2200 40.8150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.6150 73.2200 39.9150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.4160 73.2200 41.7150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.2150 73.2200 43.5160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.3150 73.2200 42.6160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.7160 73.2200 48.0170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.1150 73.2200 44.4150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.8150 73.2200 47.1140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.0150 73.2200 45.3150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.9160 73.2200 46.2160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.6150 73.2200 48.9150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.5150 73.2200 49.8150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.4160 73.2200 50.7160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.3150 73.2200 51.6140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.1150 73.2200 53.4150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.2160 73.2200 52.5170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.6150 73.2200 57.9150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.8150 73.2200 56.1140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.0150 73.2200 54.3150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.9160 73.2200 55.2160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.7150 73.2200 57.0150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.5160 73.2200 58.8160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.1150 73.2200 62.4150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.4150 73.2200 59.7140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.2150 73.2200 61.5150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.0160 73.2200 63.3160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.3160 73.2200 60.6170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.6160 73.2200 66.9160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.9150 73.2200 64.2140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.5150 73.2200 67.8140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.8150 73.2200 65.1150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.7150 73.2200 66.0150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.0150 73.2200 72.3140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.2150 73.2200 70.5150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.3150 73.2200 69.6150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.1160 73.2200 71.4160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.4160 73.2200 68.7170 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.7150 73.2200 75.0150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.6140 73.2200 75.9130 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.4140 73.2200 77.7140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.5150 73.2200 76.8160 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.9140 73.2200 73.2140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.8140 73.2200 74.1140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.1140 73.2200 80.4130 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.3140 73.2200 78.6140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.2150 73.2200 79.5150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.0140 73.2200 81.3140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.9140 73.2200 82.2140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.8150 73.2200 83.1150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.4140 73.2200 86.7140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.7140 73.2200 84.0130 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.5140 73.2200 85.8140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.3150 73.2200 87.6150 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.2140 73.2200 88.5130 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.1150 73.2200 89.4140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.0150 73.2200 90.3140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.9150 73.2200 91.2140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.8150 73.2200 92.1140 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.6150 73.2200 84.9160 73.5200 ;
    END
  END VSS

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0000 51.2600 0.2000 51.4600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0000 42.6960 0.2000 42.8960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0000 50.0630 0.2000 50.2630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.1330 0.0000 34.3330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.1330 0.0000 34.3330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.1330 0.0000 34.3330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.1330 0.0000 34.3330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.1330 0.0000 34.3330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[7]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.5010 0.0000 35.7010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.5010 0.0000 35.7010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.5010 0.0000 35.7010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.5010 0.0000 35.7010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.5010 0.0000 35.7010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[5]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.0190 0.0000 35.2190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.0190 0.0000 35.2190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.0190 0.0000 35.2190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.0190 0.0000 35.2190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.0190 0.0000 35.2190 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.5470 0.0000 29.7470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.5470 0.0000 29.7470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.5470 0.0000 29.7470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.5470 0.0000 29.7470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.5470 0.0000 29.7470 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[2]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.1790 0.0000 28.3790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.1790 0.0000 28.3790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.1790 0.0000 28.3790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.1790 0.0000 28.3790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.1790 0.0000 28.3790 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[15]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.9250 0.0000 26.1250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.9250 0.0000 26.1250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.9250 0.0000 26.1250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.9250 0.0000 26.1250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.9250 0.0000 26.1250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[6]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.8110 0.0000 27.0110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.8110 0.0000 27.0110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.8110 0.0000 27.0110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.8110 0.0000 27.0110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.8110 0.0000 27.0110 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[6]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.2930 0.0010 27.4930 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.2930 0.0010 27.4930 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.2930 0.0000 27.4930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.2930 0.0000 27.4930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.2930 0.0000 27.4930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[15]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.0290 0.0000 30.2290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.0290 0.0000 30.2290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.0290 0.0000 30.2290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.0290 0.0000 30.2290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.0290 0.0000 30.2290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[4]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.4850 0.2000 32.6850 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 32.4850 0.2000 32.6850 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 32.4850 0.2000 32.6850 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.4850 0.2000 32.6850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 32.4850 0.2000 32.6850 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[4]

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 66.5120 93.4790 66.7120 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 66.5120 93.4790 66.7120 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 66.5120 93.4790 66.7120 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 66.5120 93.4790 66.7120 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 66.5120 93.4790 66.7120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 63.3240 93.4790 63.5240 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 63.3240 93.4790 63.5240 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 63.3240 93.4790 63.5240 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 63.3240 93.4790 63.5240 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 63.3240 93.4790 63.5240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 62.9840 93.4790 63.1840 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 62.9840 93.4790 63.1840 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 62.9840 93.4790 63.1840 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 62.9840 93.4790 63.1840 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 62.9840 93.4790 63.1840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 66.5270 0.2000 66.7270 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 66.5270 0.2000 66.7270 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 66.5270 0.2000 66.7270 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 66.5270 0.2000 66.7270 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 66.5270 0.2000 66.7270 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 63.3130 0.2000 63.5130 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 63.3130 0.2000 63.5130 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 63.3130 0.2000 63.5130 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 63.3130 0.2000 63.5130 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 63.3130 0.2000 63.5130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.6360 0.0000 23.8360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.6360 0.0000 23.8360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.6360 0.0000 23.8360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.6360 0.0000 23.8360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.6360 0.0000 23.8360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 9.5898 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 60.53434 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 60.53434 LAYER M2 ;
    ANTENNAMAXAREACAR 41.79569 LAYER M2 ;
    ANTENNAGATEAREA 22.3422 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 16.28746 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.28746 LAYER M3 ;
    ANTENNAMAXAREACAR 11.33819 LAYER M3 ;
    ANTENNAGATEAREA 22.3422 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 109.4161 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 109.4161 LAYER M4 ;
    ANTENNAMAXAREACAR 47.42195 LAYER M4 ;
    ANTENNAGATEAREA 44.5773 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 3274.721 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 3274.721 LAYER M5 ;
    ANTENNAMAXAREACAR 159.7793 LAYER M5 ;
    ANTENNAGATEAREA 44.5773 LAYER M6 ;
    ANTENNAGATEAREA 44.5773 LAYER M7 ;
    ANTENNAGATEAREA 44.5773 LAYER M8 ;
    ANTENNAGATEAREA 44.5773 LAYER M9 ;
    ANTENNAGATEAREA 44.5773 LAYER MRDL ;
  END WEB2

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.9630 0.0000 46.1630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.9630 0.0000 46.1630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.9630 0.0000 46.1630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.9630 0.0000 46.1630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.9630 0.0000 46.1630 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.0770 0.0000 45.2770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.0770 0.0000 45.2770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.0770 0.0000 45.2770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.0770 0.0000 45.2770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.0770 0.0000 45.2770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.2270 0.0000 43.4270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.2270 0.0000 43.4270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.2270 0.0000 43.4270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.2270 0.0000 43.4270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.2270 0.0000 43.4270 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.7090 0.0000 43.9090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.7090 0.0000 43.9090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.7090 0.0000 43.9090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.7090 0.0000 43.9090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.7090 0.0000 43.9090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.5950 0.0000 44.7950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.5950 0.0000 44.7950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.5950 0.0000 44.7950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.5950 0.0000 44.7950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.5950 0.0000 44.7950 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.7550 0.0000 37.9550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.7550 0.0000 37.9550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.7550 0.0000 37.9550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.7550 0.0000 37.9550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.7550 0.0000 37.9550 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26404 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.8690 0.0000 37.0690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.8690 0.0000 37.0690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.8690 0.0000 37.0690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.8690 0.0000 37.0690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.8690 0.0000 37.0690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.2370 0.0000 38.4370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.2370 0.0000 38.4370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.2370 0.0000 38.4370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.2370 0.0000 38.4370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.2370 0.0000 38.4370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.3870 0.0000 36.5870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.3870 0.0000 36.5870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.3870 0.0000 36.5870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.3870 0.0000 36.5870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.3870 0.0000 36.5870 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26404 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.9730 0.0000 41.1730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.9730 0.0000 41.1730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.9730 0.0000 41.1730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.9730 0.0000 41.1730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.9730 0.0000 41.1730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.4910 0.0000 40.6910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.4910 0.0000 40.6910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.4910 0.0000 40.6910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.4910 0.0000 40.6910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.4910 0.0000 40.6910 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.6050 0.0000 39.8050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.6050 0.0000 39.8050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.6050 0.0000 39.8050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.6050 0.0000 39.8050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.6050 0.0000 39.8050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.1230 0.0000 39.3230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.1230 0.0000 39.3230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.1230 0.0000 39.3230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.1230 0.0000 39.3230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.1230 0.0000 39.3230 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26404 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.2830 0.0000 32.4830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.2830 0.0000 32.4830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.2830 0.0000 32.4830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.2830 0.0000 32.4830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.2830 0.0000 32.4830 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[11]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.3970 0.0000 31.5970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.3970 0.0000 31.5970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.3970 0.0000 31.5970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.3970 0.0000 31.5970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.3970 0.0000 31.5970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.7650 0.0000 32.9650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.7650 0.0000 32.9650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.7650 0.0000 32.9650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.7650 0.0000 32.9650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.7650 0.0000 32.9650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.6510 0.0000 33.8510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.6510 0.0000 33.8510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.6510 0.0000 33.8510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.6510 0.0000 33.8510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.6510 0.0000 33.8510 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.9150 0.0000 31.1150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.9150 0.0000 31.1150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.9150 0.0000 31.1150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.9150 0.0000 31.1150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.9150 0.0000 31.1150 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[4]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.7400 0.0000 55.9400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.7400 0.0000 55.9400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.7400 0.0000 55.9400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.7400 0.0000 55.9400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.7400 0.0000 55.9400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.0550 0.0000 55.2550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.0550 0.0000 55.2550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.0550 0.0000 55.2550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.0550 0.0000 55.2550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.0550 0.0000 55.2550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.7910 0.0000 57.9910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.7910 0.0000 57.9910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.7910 0.0000 57.9910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.7910 0.0000 57.9910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.7910 0.0000 57.9910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.1080 0.0000 57.3080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.1080 0.0000 57.3080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.1080 0.0000 57.3080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.1080 0.0000 57.3080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.1080 0.0000 57.3080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.4230 0.0000 56.6230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.4230 0.0000 56.6230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.4230 0.0000 56.6230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.4230 0.0000 56.6230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.4230 0.0000 56.6230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3720 0.0000 54.5720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.3720 0.0000 54.5720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.3720 0.0000 54.5720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.3720 0.0000 54.5720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.3720 0.0000 54.5720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.6870 0.0000 53.8870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.6870 0.0000 53.8870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.6870 0.0000 53.8870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.6870 0.0000 53.8870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.6870 0.0000 53.8870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.0040 0.0000 53.2040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.0040 0.0000 53.2040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.0040 0.0000 53.2040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.0040 0.0000 53.2040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.0040 0.0000 53.2040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.9510 0.0000 51.1510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.9510 0.0000 51.1510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.9510 0.0000 51.1510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.9510 0.0000 51.1510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.9510 0.0000 51.1510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.2680 0.0000 50.4680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.2680 0.0000 50.4680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.2680 0.0000 50.4680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.2680 0.0000 50.4680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.2680 0.0000 50.4680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.5830 0.0000 49.7830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.5830 0.0000 49.7830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.5830 0.0000 49.7830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.5830 0.0000 49.7830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.5830 0.0000 49.7830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.9000 0.0000 49.1000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.9000 0.0000 49.1000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.9000 0.0000 49.1000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.9000 0.0000 49.1000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.9000 0.0000 49.1000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.2150 0.0000 48.4150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.2150 0.0000 48.4150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.2150 0.0000 48.4150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.2150 0.0000 48.4150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.2150 0.0000 48.4150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.3140 0.0000 47.5140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.3140 0.0000 47.5140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.3140 0.0000 47.5140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.3140 0.0000 47.5140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.3140 0.0000 47.5140 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.3190 0.0000 52.5190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.3190 0.0000 52.5190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.3190 0.0000 52.5190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.3190 0.0000 52.5190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.3190 0.0000 52.5190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.6360 0.0000 51.8360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.6360 0.0000 51.8360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.6360 0.0000 51.8360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.6360 0.0000 51.8360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.6360 0.0000 51.8360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.3410 0.0000 42.5410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.3410 0.0000 42.5410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.3410 0.0000 42.5410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.3410 0.0000 42.5410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.3410 0.0000 42.5410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.8590 0.0000 42.0590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.8590 0.0000 42.0590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.8590 0.0000 42.0590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.8590 0.0000 42.0590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.8590 0.0000 42.0590 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.286324 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.4450 0.0000 46.6450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.4450 0.0000 46.6450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.4450 0.0000 46.6450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.4450 0.0000 46.6450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.4450 0.0000 46.6450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.6610 0.0000 28.8610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.6610 0.0000 28.8610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.6610 0.0000 28.8610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.6610 0.0000 28.8610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.3670 0.0000 67.5670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.3670 0.0000 67.5670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.3670 0.0000 67.5670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.3670 0.0000 67.5670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.3670 0.0000 67.5670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.6840 0.0000 66.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.6840 0.0000 66.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.6840 0.0000 66.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.6840 0.0000 66.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.6840 0.0000 66.8840 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O1[8]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.7350 0.0000 68.9350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.7350 0.0000 68.9350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.7350 0.0000 68.9350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.7350 0.0000 68.9350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.7350 0.0000 68.9350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.9480 0.0000 64.1480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.9480 0.0000 64.1480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.9480 0.0000 64.1480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.9480 0.0000 64.1480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.9480 0.0000 64.1480 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O1[14]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.0520 0.0000 68.2520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.0520 0.0000 68.2520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.0520 0.0000 68.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.0520 0.0000 68.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.0520 0.0000 68.2520 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O1[10]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.9990 0.0000 66.1990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.9990 0.0000 66.1990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.9990 0.0000 66.1990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.9990 0.0000 66.1990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.9990 0.0000 66.1990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.4200 0.0000 69.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.4200 0.0000 69.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.4200 0.0000 69.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.4200 0.0000 69.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.4200 0.0000 69.6200 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O1[3]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.3160 0.0000 65.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.3160 0.0000 65.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.3160 0.0000 65.5160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.3160 0.0000 65.5160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.3160 0.0000 65.5160 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O1[9]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.6310 0.0000 64.8310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.6310 0.0000 64.8310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.6310 0.0000 64.8310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.6310 0.0000 64.8310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.6310 0.0000 64.8310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.1590 0.0000 59.3590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.1590 0.0000 59.3590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.1590 0.0000 59.3590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.1590 0.0000 59.3590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.1590 0.0000 59.3590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.2120 0.0000 61.4120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.2120 0.0000 61.4120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.2120 0.0000 61.4120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.2120 0.0000 61.4120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.2120 0.0000 61.4120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.5270 0.0000 60.7270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.5270 0.0000 60.7270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.5270 0.0000 60.7270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.5270 0.0000 60.7270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.5270 0.0000 60.7270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.8440 0.0000 60.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.8440 0.0000 60.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.8440 0.0000 60.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.8440 0.0000 60.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.8440 0.0000 60.0440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.2630 0.0000 63.4630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.2630 0.0000 63.4630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.2630 0.0000 63.4630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.2630 0.0000 63.4630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.2630 0.0000 63.4630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.5800 0.0000 62.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.5800 0.0000 62.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.5800 0.0000 62.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.5800 0.0000 62.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.5800 0.0000 62.7800 0.2000 ;
    END
    ANTENNADIFFAREA 69.68586 LAYER M3 ;
    ANTENNADIFFAREA 70.86852 LAYER M4 ;
    ANTENNADIFFAREA 70.86852 LAYER M5 ;
    ANTENNADIFFAREA 70.86852 LAYER M6 ;
    ANTENNADIFFAREA 70.86852 LAYER M7 ;
    ANTENNADIFFAREA 70.86852 LAYER M8 ;
    ANTENNADIFFAREA 70.86852 LAYER M9 ;
    ANTENNADIFFAREA 70.86852 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 22.1883 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 12.53665 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.53665 LAYER M3 ;
    ANTENNAMAXAREACAR 7.115183 LAYER M3 ;
    ANTENNAGATEAREA 22.1883 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 91.54191 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 91.54191 LAYER M4 ;
    ANTENNAMAXAREACAR 46.54153 LAYER M4 ;
    ANTENNAGATEAREA 22.1883 LAYER M5 ;
    ANTENNAGATEAREA 22.1883 LAYER M6 ;
    ANTENNAGATEAREA 22.1883 LAYER M7 ;
    ANTENNAGATEAREA 22.1883 LAYER M8 ;
    ANTENNAGATEAREA 22.1883 LAYER M9 ;
    ANTENNAGATEAREA 22.1883 LAYER MRDL ;
  END O1[0]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.4760 0.0000 58.6760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.4760 0.0000 58.6760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.4760 0.0000 58.6760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.4760 0.0000 58.6760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.4760 0.0000 58.6760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.8950 0.0000 62.0950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.8950 0.0000 62.0950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.8950 0.0000 62.0950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.8950 0.0000 62.0950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.8950 0.0000 62.0950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2790 9.8210 93.4790 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2790 9.8210 93.4790 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2790 9.8210 93.4790 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2790 9.8210 93.4790 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2790 9.8210 93.4790 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 9.4359 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 59.36605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.36605 LAYER M2 ;
    ANTENNAMAXAREACAR 41.85088 LAYER M2 ;
    ANTENNAGATEAREA 9.4359 LAYER M3 ;
    ANTENNAGATEAREA 9.4359 LAYER M4 ;
    ANTENNAGATEAREA 9.4359 LAYER M5 ;
    ANTENNAGATEAREA 9.4359 LAYER M6 ;
    ANTENNAGATEAREA 9.4359 LAYER M7 ;
    ANTENNAGATEAREA 9.4359 LAYER M8 ;
    ANTENNAGATEAREA 9.4359 LAYER M9 ;
    ANTENNAGATEAREA 9.4359 LAYER MRDL ;
  END WEB1

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 17.5640 73.2200 17.8640 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8650 73.2200 6.1650 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9630 73.2200 5.2640 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4640 73.2200 18.7640 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.6650 73.2200 88.9650 73.5200 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.5640 73.2200 89.8640 73.5200 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 130.6569 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 130.6569 LAYER M5 ;
  END VDDL

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.46786 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.46786 LAYER M4 ;
    ANTENNAMAXAREACAR 17.30994 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 21.74154 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2
  OBS
    LAYER M2 ;
      RECT 0.0000 33.3850 93.4790 41.9130 ;
      RECT 0.9000 31.7850 92.5790 33.3850 ;
      RECT 0.9000 18.2680 92.5790 33.3850 ;
      RECT 0.9000 41.9960 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 93.4790 16.1310 ;
      RECT 0.0000 0.0000 22.9360 9.1210 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.0000 0.9000 93.4790 9.1210 ;
      RECT 0.9000 9.1210 92.5790 16.1310 ;
      RECT 0.9000 9.1210 92.5790 10.7210 ;
      RECT 70.8000 0.0000 93.4790 9.1210 ;
      RECT 70.8000 0.0000 93.4790 0.9000 ;
      RECT 0.0000 43.5960 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 43.5960 ;
      RECT 0.0000 67.4270 93.4790 73.5200 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 64.2240 ;
      RECT 0.0000 52.1600 93.4790 57.7900 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 92.5790 50.3650 93.4790 50.5600 ;
      RECT 24.5360 0.0000 25.2250 0.9000 ;
      RECT 91.9780 64.2240 93.4790 65.8120 ;
      RECT 0.0000 59.3900 93.4790 62.2840 ;
      RECT 0.0000 46.3620 92.5790 49.3630 ;
      RECT 0.9000 67.4120 93.4790 70.4130 ;
      RECT 0.0000 62.2840 92.5790 62.6130 ;
      RECT 0.9000 57.7900 92.5790 59.3900 ;
      RECT 0.0000 64.2130 1.5010 65.8270 ;
      RECT 0.0000 0.0000 22.9360 0.9000 ;
      RECT 0.0000 18.2680 93.4790 31.7850 ;
      RECT 0.0000 16.1310 92.5790 16.1340 ;
      RECT 0.9000 18.1900 93.4790 18.2680 ;
      RECT 0.9000 16.1340 92.5790 18.1900 ;
      RECT 0.0000 41.9130 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
    LAYER M1 ;
      RECT 92.6790 50.2650 93.4790 50.6600 ;
      RECT 24.4360 0.0000 25.3250 0.8000 ;
      RECT 91.9780 64.1240 93.4790 65.9120 ;
      RECT 0.0000 59.7120 92.6790 62.7130 ;
      RECT 0.0000 46.4620 92.6790 49.4630 ;
      RECT 0.8000 67.3120 93.4790 70.3130 ;
      RECT 0.0000 64.1130 1.5010 65.9270 ;
      RECT 0.0000 0.0000 23.0360 0.8000 ;
      RECT 0.0000 16.2310 92.6790 16.2340 ;
      RECT 0.0000 10.6210 92.6790 16.2340 ;
      RECT 0.0000 10.6210 92.6790 16.2340 ;
      RECT 0.0000 10.6210 92.6790 16.2340 ;
      RECT 0.0000 10.6210 93.4790 16.2310 ;
      RECT 0.0000 0.0000 23.0360 9.2210 ;
      RECT 0.8000 16.2340 92.6790 18.0900 ;
      RECT 0.8000 10.6210 92.6790 18.0900 ;
      RECT 0.8000 10.6210 92.6790 18.0900 ;
      RECT 0.8000 10.6210 92.6790 18.0900 ;
      RECT 0.0000 42.0130 92.6790 42.0960 ;
      RECT 0.8000 42.0960 92.6790 43.4130 ;
      RECT 0.0000 33.2850 92.6790 42.0960 ;
      RECT 0.0000 33.2850 92.6790 42.0960 ;
      RECT 0.0000 33.2850 92.6790 42.0960 ;
      RECT 0.0000 33.2850 93.4790 42.0130 ;
      RECT 0.0000 18.1680 93.4790 31.8850 ;
      RECT 0.8000 33.2850 92.6790 43.4130 ;
      RECT 0.8000 33.2850 92.6790 43.4130 ;
      RECT 0.8000 33.2850 92.6790 43.4130 ;
      RECT 0.8000 31.8850 92.6790 33.2850 ;
      RECT 0.8000 18.1680 92.6790 33.2850 ;
      RECT 0.8000 18.0900 93.4790 18.1680 ;
      RECT 0.0000 52.0600 93.4790 57.8900 ;
      RECT 0.8000 50.2650 92.6790 57.8900 ;
      RECT 0.8000 50.2650 92.6790 57.8900 ;
      RECT 0.8000 50.2650 92.6790 57.8900 ;
      RECT 0.8000 50.2650 92.6790 57.8900 ;
      RECT 0.0000 0.8000 93.4790 9.2210 ;
      RECT 0.8000 9.2210 92.6790 16.2310 ;
      RECT 0.8000 9.2210 92.6790 10.6210 ;
      RECT 70.7000 0.0000 93.4790 9.2210 ;
      RECT 70.7000 0.0000 93.4790 0.8000 ;
      RECT 0.0000 43.4960 93.4790 48.8650 ;
      RECT 0.8000 49.4630 92.6790 57.8900 ;
      RECT 0.8000 49.4630 92.6790 57.8900 ;
      RECT 0.8000 49.4630 92.6790 57.8900 ;
      RECT 0.8000 49.4630 92.6790 57.8900 ;
      RECT 0.8000 43.4130 93.4790 48.8650 ;
      RECT 0.8000 43.4130 93.4790 48.8650 ;
      RECT 0.8000 43.4130 93.4790 48.8650 ;
      RECT 0.8000 43.4130 93.4790 43.4960 ;
      RECT 0.0000 67.3270 93.4790 73.5200 ;
      RECT 0.0000 59.2900 93.4790 62.3840 ;
      RECT 0.8000 64.1130 92.6790 67.3120 ;
      RECT 0.8000 64.1130 92.6790 67.3120 ;
      RECT 0.8000 64.1130 92.6790 67.3120 ;
      RECT 0.8000 64.1130 92.6790 67.3120 ;
      RECT 0.8000 64.1130 92.6790 67.3120 ;
      RECT 0.8000 62.7130 92.6790 67.3120 ;
      RECT 0.8000 62.7130 92.6790 67.3120 ;
      RECT 0.8000 62.7130 92.6790 67.3120 ;
      RECT 0.8000 62.7130 92.6790 67.3120 ;
      RECT 0.8000 62.7130 92.6790 67.3120 ;
      RECT 0.8000 64.1130 92.6790 64.1240 ;
      RECT 0.8000 57.8900 92.6790 62.3840 ;
      RECT 0.8000 57.8900 92.6790 59.2900 ;
    LAYER PO ;
      RECT 0.0000 0.0000 93.4790 73.5200 ;
    LAYER M4 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 93.4790 16.1310 ;
      RECT 0.9000 18.1900 93.4790 18.2680 ;
      RECT 0.9000 16.1340 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.0000 0.9010 93.4790 9.1210 ;
      RECT 0.9000 9.1210 92.5790 16.1310 ;
      RECT 0.9000 9.1210 92.5790 10.7210 ;
      RECT 28.1930 0.9000 93.4790 9.1210 ;
      RECT 28.1930 0.9000 93.4790 9.1210 ;
      RECT 28.1930 0.9000 93.4790 9.1210 ;
      RECT 28.1930 0.9000 93.4790 0.9010 ;
      RECT 70.8000 0.0000 93.4790 9.1210 ;
      RECT 70.8000 0.0000 93.4790 9.1210 ;
      RECT 70.8000 0.0000 93.4790 0.9000 ;
      RECT 0.9000 64.2240 92.5790 65.8120 ;
      RECT 0.0000 43.5960 93.4790 48.7650 ;
      RECT 0.9000 50.3650 92.5790 50.5600 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 43.5960 ;
      RECT 0.9000 65.8120 92.5790 65.8270 ;
      RECT 0.9000 64.2130 92.5790 64.2240 ;
      RECT 0.0000 67.4270 93.4790 73.5200 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.0000 52.1600 93.4790 57.7900 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 24.5360 0.0000 25.2250 0.9000 ;
      RECT 0.0000 62.2840 92.5790 62.6130 ;
      RECT 0.0000 46.3620 92.5790 49.3630 ;
      RECT 0.0000 59.3900 93.4790 62.2840 ;
      RECT 0.0000 64.2130 1.5010 65.8270 ;
      RECT 0.9000 50.3650 93.4790 50.5600 ;
      RECT 0.9000 49.3630 92.5790 50.3650 ;
      RECT 0.9000 57.7900 92.5790 59.3900 ;
      RECT 0.9000 67.4120 93.4790 70.4130 ;
      RECT 0.9000 50.5600 92.5790 50.8640 ;
      RECT 91.9780 64.2240 93.4790 65.8120 ;
      RECT 0.0000 0.0000 22.9360 0.9000 ;
      RECT 0.0000 0.9000 26.5930 0.9010 ;
      RECT 0.0000 0.0000 22.9360 9.1210 ;
      RECT 0.0000 0.0000 22.9360 9.1210 ;
      RECT 0.0000 0.9000 26.5930 9.1210 ;
      RECT 0.0000 0.9000 26.5930 9.1210 ;
      RECT 0.0000 0.9000 26.5930 9.1210 ;
      RECT 0.0000 18.2680 93.4790 31.7850 ;
      RECT 0.0000 41.9130 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 93.4790 41.9130 ;
      RECT 0.9000 41.9960 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 31.7850 92.5790 41.9130 ;
      RECT 0.9000 31.7850 92.5790 33.3850 ;
      RECT 0.0000 16.1310 92.5790 16.1340 ;
    LAYER M3 ;
      RECT 24.5360 0.0000 25.2250 0.9000 ;
      RECT 0.0000 62.2840 92.5790 62.6130 ;
      RECT 0.0000 46.3620 92.5790 49.3630 ;
      RECT 0.0000 59.3900 93.4790 62.2840 ;
      RECT 0.0000 64.2130 1.5010 65.8270 ;
      RECT 0.9000 57.7900 92.5790 59.3900 ;
      RECT 0.9000 67.4120 93.4790 70.4130 ;
      RECT 91.9780 64.2240 93.4790 65.8120 ;
      RECT 92.5790 50.3650 93.4790 50.5600 ;
      RECT 0.0000 0.0000 22.9360 0.9000 ;
      RECT 0.0000 18.2680 93.4790 31.7850 ;
      RECT 0.0000 16.1310 92.5790 16.1340 ;
      RECT 0.9000 18.1900 93.4790 18.2680 ;
      RECT 0.9000 16.1340 92.5790 18.1900 ;
      RECT 0.0000 41.9130 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 93.4790 41.9130 ;
      RECT 0.9000 31.7850 92.5790 33.3850 ;
      RECT 0.9000 18.2680 92.5790 33.3850 ;
      RECT 0.9000 41.9960 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 93.4790 16.1310 ;
      RECT 0.0000 0.0000 22.9360 9.1210 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.0000 0.9000 93.4790 9.1210 ;
      RECT 0.9000 9.1210 92.5790 16.1310 ;
      RECT 0.9000 9.1210 92.5790 10.7210 ;
      RECT 70.8000 0.0000 93.4790 9.1210 ;
      RECT 70.8000 0.0000 93.4790 0.9000 ;
      RECT 0.0000 43.5960 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 43.5960 ;
      RECT 0.0000 67.4270 93.4790 73.5200 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 67.4120 ;
      RECT 0.9000 64.2130 92.5790 64.2240 ;
      RECT 0.0000 52.1600 93.4790 57.7900 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
      RECT 0.9000 49.3630 92.5790 57.7900 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 93.4790 73.5200 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 93.4790 73.5200 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 93.4790 73.5200 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 93.4790 73.5200 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 93.4790 73.5200 ;
    LAYER M5 ;
      RECT 93.2650 72.5200 93.4790 73.5200 ;
      RECT 0.0000 72.5200 0.6630 73.5200 ;
      RECT 24.5360 0.0000 25.2250 0.9000 ;
      RECT 0.0000 59.3900 3.0010 62.6130 ;
      RECT 0.0000 46.3620 92.5790 49.3630 ;
      RECT 0.0000 64.2130 1.5010 65.8270 ;
      RECT 0.9000 50.3650 93.4790 50.5600 ;
      RECT 0.9000 49.3630 92.5790 50.3650 ;
      RECT 0.9000 67.4120 93.4790 70.4130 ;
      RECT 0.9000 50.5600 92.5790 50.8640 ;
      RECT 91.9780 64.2240 93.4790 65.8120 ;
      RECT 91.9780 59.3900 93.4790 62.2840 ;
      RECT 0.0000 0.9000 26.5930 0.9010 ;
      RECT 0.0000 0.0000 22.9360 0.9000 ;
      RECT 0.0000 18.2680 93.4790 31.7850 ;
      RECT 0.9000 18.1900 93.4790 18.2680 ;
      RECT 0.9000 16.1340 92.5790 18.1900 ;
      RECT 0.0000 16.1310 92.5790 16.1340 ;
      RECT 0.0000 41.9130 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 92.5790 41.9960 ;
      RECT 0.0000 33.3850 93.4790 41.9130 ;
      RECT 0.9000 31.7850 92.5790 41.9130 ;
      RECT 0.9000 31.7850 92.5790 33.3850 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 92.5790 16.1340 ;
      RECT 0.0000 10.7210 93.4790 16.1310 ;
      RECT 0.0000 0.0000 22.9360 9.1210 ;
      RECT 0.0000 0.0000 22.9360 9.1210 ;
      RECT 0.0000 0.9000 26.5930 9.1210 ;
      RECT 0.0000 0.9000 26.5930 9.1210 ;
      RECT 0.0000 0.9000 26.5930 9.1210 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 10.7210 92.5790 18.1900 ;
      RECT 0.9000 41.9960 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.9000 33.3850 92.5790 43.5130 ;
      RECT 0.0000 0.9010 93.4790 9.1210 ;
      RECT 0.9000 9.1210 92.5790 16.1310 ;
      RECT 0.9000 9.1210 92.5790 10.7210 ;
      RECT 28.1930 0.9000 93.4790 9.1210 ;
      RECT 28.1930 0.9000 93.4790 9.1210 ;
      RECT 28.1930 0.9000 93.4790 9.1210 ;
      RECT 28.1930 0.9000 93.4790 0.9010 ;
      RECT 70.8000 0.0000 93.4790 9.1210 ;
      RECT 70.8000 0.0000 93.4790 9.1210 ;
      RECT 70.8000 0.0000 93.4790 0.9000 ;
      RECT 0.9000 64.2240 92.5790 65.8120 ;
      RECT 0.9000 64.2130 92.5790 64.2240 ;
      RECT 0.9000 62.6130 92.5790 65.8120 ;
      RECT 0.9000 62.6130 92.5790 65.8120 ;
      RECT 0.9000 62.2840 92.5790 65.8120 ;
      RECT 0.9000 62.2840 92.5790 65.8120 ;
      RECT 0.9000 62.2840 92.5790 65.8120 ;
      RECT 0.9000 62.2840 92.5790 65.8120 ;
      RECT 0.0000 43.5960 93.4790 48.7650 ;
      RECT 0.9000 50.3650 92.5790 50.5600 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 48.7650 ;
      RECT 0.9000 43.5130 93.4790 43.5960 ;
      RECT 0.0000 67.4270 93.4790 72.5200 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 64.2240 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.9000 62.6130 92.5790 67.4120 ;
      RECT 0.0000 52.1600 93.4790 57.7900 ;
      RECT 0.9000 59.3900 92.5790 65.8120 ;
      RECT 0.9000 57.7900 92.5790 65.8120 ;
      RECT 0.9000 57.7900 92.5790 65.8120 ;
      RECT 0.9000 57.7900 92.5790 62.2840 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
      RECT 0.9000 50.3650 92.5790 57.7900 ;
  END
END SRAMLP2RW32x16

MACRO SRAMLP2RW32x22
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 104.046 BY 74.598 ;
  SYMMETRY X Y R90 ;

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[14]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.4700 0.0000 57.6700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.4700 0.0000 57.6700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.4700 0.0000 57.6700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.4700 0.0000 57.6700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.4700 0.0000 57.6700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[21]

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.2600 0.0020 83.4600 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.2600 0.0020 83.4600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.2600 0.0020 83.4600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.2600 0.0020 83.4600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.2600 0.0020 83.4600 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.3618 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.0605 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0605 LAYER M2 ;
    ANTENNAMAXAREACAR 6.661157 LAYER M2 ;
    ANTENNAGATEAREA 0.3618 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 7.079733 LAYER M3 ;
    ANTENNAGATEAREA 0.3618 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.498282 LAYER M4 ;
    ANTENNAGATEAREA 0.3618 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.916803 LAYER M5 ;
    ANTENNAGATEAREA 0.3618 LAYER M6 ;
    ANTENNAGATEAREA 0.3618 LAYER M7 ;
    ANTENNAGATEAREA 0.3618 LAYER M8 ;
    ANTENNAGATEAREA 0.3618 LAYER M9 ;
    ANTENNAGATEAREA 0.3618 LAYER MRDL ;
  END OEB1

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5800 0.0020 20.7800 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5800 0.0020 20.7800 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5800 0.0020 20.7800 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5800 0.0020 20.7800 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5800 0.0020 20.7800 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.3618 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.06026 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.06026 LAYER M2 ;
    ANTENNAMAXAREACAR 6.660493 LAYER M2 ;
    ANTENNAGATEAREA 0.3618 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 7.07907 LAYER M3 ;
    ANTENNAGATEAREA 0.3618 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.497619 LAYER M4 ;
    ANTENNAGATEAREA 0.3618 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.91614 LAYER M5 ;
    ANTENNAGATEAREA 0.3618 LAYER M6 ;
    ANTENNAGATEAREA 0.3618 LAYER M7 ;
    ANTENNAGATEAREA 0.3618 LAYER M8 ;
    ANTENNAGATEAREA 0.3618 LAYER M9 ;
    ANTENNAGATEAREA 0.3618 LAYER MRDL ;
  END OEB2

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 9.8950 104.0460 10.0950 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 9.8950 104.0460 10.0950 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 9.8950 104.0460 10.0950 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 9.8950 104.0460 10.0950 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 9.8950 104.0460 10.0950 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16072 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16072 LAYER M1 ;
    ANTENNAGATEAREA 0.1704 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.60152 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.60152 LAYER M2 ;
    ANTENNAMAXAREACAR 11.94964 LAYER M2 ;
    ANTENNAGATEAREA 0.1704 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.15352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15352 LAYER M3 ;
    ANTENNAMAXAREACAR 12.8498 LAYER M3 ;
    ANTENNAGATEAREA 0.1704 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.15352 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15352 LAYER M4 ;
    ANTENNAMAXAREACAR 13.74991 LAYER M4 ;
    ANTENNAGATEAREA 0.1704 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.15352 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15352 LAYER M5 ;
    ANTENNAMAXAREACAR 14.64995 LAYER M5 ;
    ANTENNAGATEAREA 0.1704 LAYER M6 ;
    ANTENNAGATEAREA 0.1704 LAYER M7 ;
    ANTENNAGATEAREA 0.1704 LAYER M8 ;
    ANTENNAGATEAREA 0.1704 LAYER M9 ;
    ANTENNAGATEAREA 0.1704 LAYER MRDL ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAGATEAREA 0.1704 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.60152 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.60152 LAYER M2 ;
    ANTENNAMAXAREACAR 11.94964 LAYER M2 ;
    ANTENNAGATEAREA 0.1704 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.83853 LAYER M3 ;
    ANTENNAGATEAREA 0.1704 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.72735 LAYER M4 ;
    ANTENNAGATEAREA 0.1704 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.61612 LAYER M5 ;
    ANTENNAGATEAREA 0.1704 LAYER M6 ;
    ANTENNAGATEAREA 0.1704 LAYER M7 ;
    ANTENNAGATEAREA 0.1704 LAYER M8 ;
    ANTENNAGATEAREA 0.1704 LAYER M9 ;
    ANTENNAGATEAREA 0.1704 LAYER MRDL ;
  END WEB2

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 54.5600 0.2000 54.7600 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 54.5600 0.2000 54.7600 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 54.5600 0.2000 54.7600 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 54.5600 0.2000 54.7600 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 54.5600 0.2000 54.7600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
  END A2[1]

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 64.7020 0.2000 64.9020 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 64.7020 0.2000 64.9020 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 64.7020 0.2000 64.9020 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 64.7020 0.2000 64.9020 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 64.7020 0.2000 64.9020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.299628 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.299628 LAYER M2 ;
    ANTENNAMAXAREACAR 15.99411 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.176024 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.176024 LAYER M3 ;
    ANTENNAMAXAREACAR 28.08656 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 45.10579 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 48.42737 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS2

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 67.9160 0.2000 68.1160 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 67.9160 0.2000 68.1160 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 67.9160 0.2000 68.1160 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 67.9160 0.2000 68.1160 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 67.9160 0.2000 68.1160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.288165 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288165 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 29.82637 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 32.86858 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.91059 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 67.9190 104.0460 68.1190 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 67.9190 104.0460 68.1190 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 67.9190 104.0460 68.1190 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 67.9190 104.0460 68.1190 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 67.9190 104.0460 68.1190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.343545 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.343545 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 31.33937 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 34.38148 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 37.42339 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 64.3650 104.0460 64.5650 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 64.3650 104.0460 64.5650 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 64.3650 104.0460 64.5650 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 64.3650 104.0460 64.5650 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 64.3650 104.0460 64.5650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.2043 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.480391 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.480391 LAYER M2 ;
    ANTENNAMAXAREACAR 9.566273 LAYER M2 ;
    ANTENNAGATEAREA 0.6282 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 6.059947 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.059947 LAYER M3 ;
    ANTENNAMAXAREACAR 17.54282 LAYER M3 ;
    ANTENNAGATEAREA 0.6282 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 19.45284 LAYER M4 ;
    ANTENNAGATEAREA 0.6282 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 19.69288 LAYER M5 ;
    ANTENNAGATEAREA 0.6282 LAYER M6 ;
    ANTENNAGATEAREA 0.6282 LAYER M7 ;
    ANTENNAGATEAREA 0.6282 LAYER M8 ;
    ANTENNAGATEAREA 0.6282 LAYER M9 ;
    ANTENNAGATEAREA 0.6282 LAYER MRDL ;
  END SD

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[20]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[19]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 35.7940 104.0460 35.9940 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 35.7940 104.0460 35.9940 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 35.7940 104.0460 35.9940 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 35.7940 104.0460 35.9940 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 35.7940 104.0460 35.9940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.08982 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.08982 LAYER M4 ;
    ANTENNAMAXAREACAR 65.87479 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 73.08949 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[4]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 61.8230 104.0460 62.0230 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 61.8230 104.0460 62.0230 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 61.8230 104.0460 62.0230 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 61.8230 104.0460 62.0230 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 61.8230 104.0460 62.0230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M2 ;
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 54.5230 104.0460 54.7230 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 54.5230 104.0460 54.7230 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 54.5230 104.0460 54.7230 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 54.5230 104.0460 54.7230 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 54.5230 104.0460 54.7230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M2 ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 52.9970 104.0460 53.1970 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 52.9970 104.0460 53.1970 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 52.9970 104.0460 53.1970 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 52.9970 104.0460 53.1970 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 52.9970 104.0460 53.1970 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M2 ;
  END A1[2]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.40684 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40684 LAYER M4 ;
    ANTENNAMAXAREACAR 13.56469 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.70587 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4090 0.2000 17.6090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4090 0.2000 17.6090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4090 0.2000 17.6090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4090 0.2000 17.6090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4090 0.2000 17.6090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30916 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30916 LAYER M4 ;
    ANTENNAMAXAREACAR 13.1427 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.57459 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 35.7540 0.2000 35.9540 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 35.7540 0.2000 35.9540 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 35.7540 0.2000 35.9540 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 35.7540 0.2000 35.9540 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 35.7540 0.2000 35.9540 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.0906 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0906 LAYER M4 ;
    ANTENNAMAXAREACAR 65.17186 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 72.3866 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[4]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 45.7350 0.2000 45.9350 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 45.7350 0.2000 45.9350 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 45.7350 0.2000 45.9350 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 45.7350 0.2000 45.9350 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 45.7350 0.2000 45.9350 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 31.9104 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 49.16678 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.16678 LAYER M3 ;
    ANTENNAMAXAREACAR 23.18403 LAYER M3 ;
    ANTENNAGATEAREA 31.9104 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 330.3812 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 330.3812 LAYER M4 ;
    ANTENNAMAXAREACAR 33.53744 LAYER M4 ;
    ANTENNAGATEAREA 40.503 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 4256.356 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 4256.356 LAYER M5 ;
    ANTENNAMAXAREACAR 192.0611 LAYER M5 ;
    ANTENNAGATEAREA 40.503 LAYER M6 ;
    ANTENNAGATEAREA 40.503 LAYER M7 ;
    ANTENNAGATEAREA 40.503 LAYER M8 ;
    ANTENNAGATEAREA 40.503 LAYER M9 ;
    ANTENNAGATEAREA 40.503 LAYER MRDL ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 53.0400 0.2000 53.2400 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 53.0400 0.2000 53.2400 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 53.0400 0.2000 53.2400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 53.0400 0.2000 53.2400 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 53.0400 0.2000 53.2400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
  END A2[2]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 61.8120 0.2000 62.0120 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 61.8120 0.2000 62.0120 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 61.8120 0.2000 62.0120 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 61.8120 0.2000 62.0120 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 61.8120 0.2000 62.0120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
  END A2[0]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 45.6960 104.0460 45.8960 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 45.6960 104.0460 45.8960 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 45.6960 104.0460 45.8960 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 45.6960 104.0460 45.8960 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 45.6960 104.0460 45.8960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M2 ;
  END A1[3]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.3660 0.0000 53.5660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.3660 0.0000 53.5660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.3660 0.0000 53.5660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.3660 0.0000 53.5660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.3660 0.0000 53.5660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[18]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 17.3650 104.0460 17.5650 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 17.3650 104.0460 17.5650 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 17.3650 104.0460 17.5650 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 17.3650 104.0460 17.5650 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 17.3650 104.0460 17.5650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.29968 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.29968 LAYER M4 ;
    ANTENNAMAXAREACAR 13.19096 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.62284 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 16.9030 104.0460 17.1030 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 16.9030 104.0460 17.1030 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 16.9030 104.0460 17.1030 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 16.9030 104.0460 17.1030 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 16.9030 104.0460 17.1030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.424789 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.424789 LAYER M4 ;
    ANTENNAMAXAREACAR 14.05956 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.20071 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 100.0070 74.2980 100.3060 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.9080 74.2980 101.2070 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8090 74.2980 12.1080 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.7090 74.2980 13.0080 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9090 74.2980 2.2080 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.8080 74.2980 3.1090 74.5980 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 5.0580 74.2980 5.3590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.1580 74.2980 4.4590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2580 74.2980 3.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3590 74.2980 2.6590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4580 74.2980 1.7580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5580 74.2980 9.8590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6580 74.2980 8.9590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4590 74.2980 10.7590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7590 74.2980 8.0580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8590 74.2980 7.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9590 74.2980 6.2590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3590 74.2980 11.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9590 74.2980 15.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0580 74.2980 14.3580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1590 74.2980 13.4590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2580 74.2980 12.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3590 74.2980 20.6590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5580 74.2980 18.8590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6580 74.2980 17.9590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7580 74.2980 17.0590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8580 74.2980 16.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4590 74.2980 19.7590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2580 74.2980 21.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8580 74.2980 25.1590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1580 74.2980 22.4590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9590 74.2980 24.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0590 74.2980 23.3590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7580 74.2980 26.0580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6590 74.2980 26.9590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5580 74.2980 27.8580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4590 74.2980 28.7590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3590 74.2980 29.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8590 74.2980 34.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9590 74.2980 33.2590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1580 74.2980 31.4590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7590 74.2980 35.0580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2590 74.2980 30.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0580 74.2980 32.3590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4580 74.2980 37.7580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6580 74.2980 35.9590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5580 74.2980 36.8590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3580 74.2980 38.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2590 74.2980 39.5590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8580 74.2980 43.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7590 74.2980 44.0590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1580 74.2980 40.4570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9580 74.2980 42.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0590 74.2980 41.3600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3580 74.2980 47.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1580 74.2980 49.4570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2590 74.2980 48.5590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4580 74.2980 46.7580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5590 74.2980 45.8600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6580 74.2980 44.9570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7590 74.2980 53.0590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9580 74.2980 51.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6580 74.2980 53.9580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8580 74.2980 52.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0590 74.2980 50.3600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0580 74.2980 59.3580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1580 74.2980 58.4580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2580 74.2980 57.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4580 74.2980 55.7580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5580 74.2980 54.8580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3590 74.2980 56.6590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6570 74.2980 62.9570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7580 74.2980 62.0580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8580 74.2980 61.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5580 74.2980 63.8580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9590 74.2980 60.2590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0590 74.2980 68.3590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1580 74.2980 67.4580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2580 74.2980 66.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3570 74.2980 65.6570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4570 74.2980 64.7570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4590 74.2980 73.7590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5580 74.2980 72.8580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6600 74.2980 71.9600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7590 74.2980 71.0590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8590 74.2980 70.1590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9580 74.2980 69.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9580 74.2980 78.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.0600 74.2980 77.3600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1590 74.2980 76.4590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2590 74.2980 75.5590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3580 74.2980 74.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4600 74.2980 82.7600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5590 74.2980 81.8590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6600 74.2980 80.9600 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7590 74.2980 80.0590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8590 74.2980 79.1590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.8570 74.2980 88.1570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.9580 74.2980 87.2580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0570 74.2980 86.3570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1580 74.2980 85.4580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2580 74.2980 84.5580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3590 74.2980 83.6590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.3580 74.2980 92.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.4570 74.2980 91.7570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.5580 74.2980 90.8580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.6570 74.2980 89.9570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.7580 74.2980 89.0580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.8580 74.2980 97.1580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.9590 74.2980 96.2590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.0570 74.2980 95.3570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.1580 74.2980 94.4580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.7590 74.2980 98.0590 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.6580 74.2980 98.9580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.5580 74.2980 99.8580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.4570 74.2980 100.7570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.3580 74.2980 101.6580 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.2570 74.2980 102.5570 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.2570 74.2980 93.5570 74.5980 ;
    END
  END VSS

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[19]

  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[17]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.9680 0.0020 65.1680 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.9680 0.0020 65.1680 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.9680 0.0020 65.1680 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.9680 0.0020 65.1680 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.9680 0.0020 65.1680 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[20]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[17]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[17]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[15]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.3360 0.0020 66.5360 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.3360 0.0020 66.5360 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.3360 0.0020 66.5360 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.3360 0.0020 66.5360 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.3360 0.0020 66.5360 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[16]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[8]

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 93.7080 74.2980 94.0070 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.6070 74.2980 94.9060 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.3090 74.2980 16.6090 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.2090 74.2980 17.5080 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.5090 74.2980 5.8080 74.5980 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.4080 74.2980 6.7090 74.5980 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 132.4626 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 132.4626 LAYER M5 ;
  END VDDL

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[11]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[18]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.1020 0.0000 56.3020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.1020 0.0000 56.3020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.1020 0.0000 56.3020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.1020 0.0000 56.3020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.1020 0.0000 56.3020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[16]

  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[21]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.0240 0.0020 54.2240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.0240 0.0020 54.2240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.0240 0.0020 54.2240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.0240 0.0020 54.2240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.0240 0.0020 54.2240 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[18]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.8460 64.7050 104.0460 64.9050 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.8460 64.7050 104.0460 64.9050 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8460 64.7050 104.0460 64.9050 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8460 64.7050 104.0460 64.9050 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8460 64.7050 104.0460 64.9050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.355008 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.355008 LAYER M2 ;
    ANTENNAMAXAREACAR 18.59413 LAYER M2 ;
    ANTENNAGATEAREA 0.132 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 5.795813 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.795813 LAYER M3 ;
    ANTENNAMAXAREACAR 56.59697 LAYER M3 ;
    ANTENNAGATEAREA 0.132 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 30.4315 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.4315 LAYER M4 ;
    ANTENNAMAXAREACAR 293.0434 LAYER M4 ;
    ANTENNAGATEAREA 0.132 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 132.6142 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 132.6142 LAYER M5 ;
    ANTENNAMAXAREACAR 1297.696 LAYER M5 ;
    ANTENNAGATEAREA 0.132 LAYER M6 ;
    ANTENNAGATEAREA 0.132 LAYER M7 ;
    ANTENNAGATEAREA 0.132 LAYER M8 ;
    ANTENNAGATEAREA 0.132 LAYER M9 ;
    ANTENNAGATEAREA 0.132 LAYER MRDL ;
  END DS1

  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.6560 0.0020 52.8560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.6560 0.0020 52.8560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.6560 0.0020 52.8560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.6560 0.0020 52.8560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.6560 0.0020 52.8560 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.301848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.301848 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[19]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[15]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[19]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.1280 0.0020 58.3280 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.1280 0.0020 58.3280 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.1280 0.0020 58.3280 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.1280 0.0020 58.3280 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.1280 0.0020 58.3280 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[21]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[17]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.6000 0.0020 63.8000 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.6000 0.0020 63.8000 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.6000 0.0020 63.8000 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.6000 0.0020 63.8000 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.6000 0.0020 63.8000 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[16]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.6780 0.0000 65.8780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.6780 0.0000 65.8780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.6780 0.0000 65.8780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.6780 0.0000 65.8780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6780 0.0000 65.8780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.2320 0.0020 62.4320 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.2320 0.0020 62.4320 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.2320 0.0020 62.4320 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.2320 0.0020 62.4320 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.2320 0.0020 62.4320 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[9]

  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[18]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.3100 0.0000 64.5100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.3100 0.0000 64.5100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.3100 0.0000 64.5100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.3100 0.0000 64.5100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.3100 0.0000 64.5100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[20]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.5740 0.0000 61.7740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.5740 0.0000 61.7740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.5740 0.0000 61.7740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.5740 0.0000 61.7740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.5740 0.0000 61.7740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[21]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.7600 0.0020 56.9600 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.7600 0.0020 56.9600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.7600 0.0020 56.9600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.7600 0.0020 56.9600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.7600 0.0020 56.9600 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[16]

  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[20]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[10]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.4960 0.0020 59.6960 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.4960 0.0020 59.6960 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.4960 0.0020 59.6960 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.4960 0.0020 59.6960 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.4960 0.0020 59.6960 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.3920 0.0020 55.5920 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.3920 0.0020 55.5920 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.3920 0.0020 55.5920 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.3920 0.0020 55.5920 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.3920 0.0020 55.5920 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.8380 0.0000 59.0380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.8380 0.0000 59.0380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.8380 0.0000 59.0380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.8380 0.0000 59.0380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.8380 0.0000 59.0380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.65304 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.65304 LAYER M3 ;
    ANTENNAMAXAREACAR 79.96445 LAYER M3 ;
    ANTENNAGATEAREA 0.4062 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 15.47993 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.47993 LAYER M4 ;
    ANTENNAMAXAREACAR 51.3611 LAYER M4 ;
    ANTENNAGATEAREA 0.4062 LAYER M5 ;
    ANTENNAGATEAREA 0.4062 LAYER M6 ;
    ANTENNAGATEAREA 0.4062 LAYER M7 ;
    ANTENNAGATEAREA 0.4062 LAYER M8 ;
    ANTENNAGATEAREA 0.4062 LAYER M9 ;
    ANTENNAGATEAREA 0.4062 LAYER MRDL ;
  END I1[1]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.2060 0.0000 60.4060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.2060 0.0000 60.4060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.2060 0.0000 60.4060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.2060 0.0000 60.4060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.2060 0.0000 60.4060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.8640 0.0020 61.0640 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.8640 0.0020 61.0640 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.8640 0.0020 61.0640 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.8640 0.0020 61.0640 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.8640 0.0020 61.0640 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7340 0.0000 54.9340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7340 0.0000 54.9340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7340 0.0000 54.9340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7340 0.0000 54.9340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7340 0.0000 54.9340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.9420 0.0000 63.1420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.9420 0.0000 63.1420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.9420 0.0000 63.1420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.9420 0.0000 63.1420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.9420 0.0000 63.1420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]
  OBS
    LAYER M2 ;
      RECT 0.9000 65.6050 103.1460 68.8190 ;
      RECT 0.9000 64.0020 103.1460 68.8190 ;
      RECT 0.9000 64.0020 103.1460 68.8190 ;
      RECT 0.9000 61.1230 103.1460 68.8190 ;
      RECT 0.9000 65.6050 103.1460 68.8160 ;
      RECT 0.9000 65.6050 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 61.1230 103.1460 67.2190 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 51.7860 0.9000 51.9560 0.9020 ;
      RECT 0.0000 62.7120 0.9000 64.0020 ;
      RECT 0.0000 68.8160 3.0010 68.8190 ;
      RECT 0.0000 65.6020 1.5010 67.2160 ;
      RECT 21.4800 0.0000 22.1680 0.9020 ;
      RECT 51.7860 0.9000 51.9560 1.0510 ;
      RECT 101.0450 61.1120 104.0460 61.1230 ;
      RECT 102.5450 65.6050 104.0460 67.2190 ;
      RECT 103.1460 62.7230 104.0460 63.6650 ;
      RECT 0.0000 52.2970 103.1460 52.3400 ;
      RECT 0.9000 35.0940 103.1460 36.6540 ;
      RECT 0.0000 44.9960 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 104.0460 44.9960 ;
      RECT 0.0000 36.6540 103.1460 36.6940 ;
      RECT 0.0000 46.6350 103.1460 52.3400 ;
      RECT 0.0000 46.6350 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 46.6350 ;
      RECT 0.9000 45.0350 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.0000 16.2030 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 104.0460 16.2030 ;
      RECT 0.0000 0.0000 19.8800 9.1950 ;
      RECT 0.0000 0.0000 19.8800 0.9020 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 10.7960 ;
      RECT 0.9000 9.1960 103.1460 10.7950 ;
      RECT 0.9000 52.3400 103.1460 55.4230 ;
      RECT 0.9000 46.6350 103.1460 55.4230 ;
      RECT 0.0000 18.3090 104.0460 35.0540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 35.0540 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 18.3090 ;
      RECT 0.9000 16.2090 103.1460 18.2650 ;
      RECT 0.0000 9.1950 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 104.0460 9.1950 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 84.1600 0.0000 104.0460 9.1950 ;
      RECT 84.1600 0.0000 104.0460 0.9020 ;
      RECT 0.0000 68.8190 104.0460 74.5980 ;
      RECT 0.0000 55.4600 104.0460 61.1120 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4230 104.0460 55.4600 ;
      RECT 0.9000 52.3400 103.1460 55.4600 ;
      RECT 0.9000 64.0020 103.1460 74.5980 ;
      RECT 0.9000 64.0020 103.1460 74.5980 ;
      RECT 0.9000 61.1230 103.1460 74.5980 ;
    LAYER M1 ;
      RECT 51.6860 0.8000 52.0560 0.8020 ;
      RECT 0.0000 68.7160 3.0010 68.7190 ;
      RECT 0.0000 53.8400 104.0460 53.9230 ;
      RECT 0.0000 53.9230 103.2460 53.9600 ;
      RECT 0.0000 52.3970 3.0010 52.4400 ;
      RECT 0.0000 62.6120 0.8000 64.1020 ;
      RECT 0.0000 65.5020 1.5010 67.3160 ;
      RECT 0.8000 53.8220 104.0460 53.8400 ;
      RECT 0.8000 53.9600 103.2460 55.3230 ;
      RECT 0.8000 55.3230 104.0460 58.3240 ;
      RECT 21.3800 0.0000 22.2680 0.8020 ;
      RECT 51.6860 0.8000 52.0560 1.1010 ;
      RECT 101.0450 61.2120 104.0460 61.2230 ;
      RECT 102.5450 65.5050 104.0460 67.3190 ;
      RECT 103.2460 62.6230 104.0460 63.7650 ;
      RECT 103.2460 53.7970 104.0460 53.8220 ;
      RECT 0.0000 36.5940 104.0460 45.0960 ;
      RECT 0.0000 45.0960 103.2460 45.1350 ;
      RECT 0.0000 36.5940 103.2460 45.1350 ;
      RECT 0.0000 36.5940 103.2460 45.1350 ;
      RECT 0.0000 36.5940 103.2460 45.1350 ;
      RECT 0.8000 53.8400 103.2460 53.9230 ;
      RECT 0.8000 53.7970 103.2460 53.8400 ;
      RECT 0.8000 45.1350 103.2460 46.4960 ;
      RECT 0.0000 36.5540 103.2460 36.5940 ;
      RECT 0.8000 16.3090 103.2460 18.1650 ;
      RECT 0.8000 18.1650 104.0460 18.2090 ;
      RECT 0.0000 16.3030 103.2460 16.3090 ;
      RECT 0.0000 10.6960 103.2460 16.3090 ;
      RECT 0.0000 10.6960 103.2460 16.3090 ;
      RECT 0.0000 10.6960 103.2460 16.3090 ;
      RECT 0.0000 10.6960 104.0460 16.3030 ;
      RECT 0.0000 0.0000 19.9800 9.2950 ;
      RECT 0.0000 0.0000 19.9800 0.8020 ;
      RECT 0.8000 10.6950 104.0460 16.3030 ;
      RECT 0.8000 10.6950 104.0460 16.3030 ;
      RECT 0.8000 10.6950 104.0460 16.3030 ;
      RECT 0.8000 10.6950 104.0460 10.6960 ;
      RECT 0.8000 9.2960 103.2460 10.6950 ;
      RECT 0.0000 18.2090 104.0460 35.1540 ;
      RECT 0.8000 35.1940 103.2460 36.5540 ;
      RECT 0.8000 18.2090 103.2460 36.5540 ;
      RECT 0.8000 18.2090 103.2460 36.5540 ;
      RECT 0.8000 18.2090 103.2460 36.5540 ;
      RECT 0.8000 35.1540 104.0460 35.1940 ;
      RECT 0.8000 18.2090 104.0460 35.1940 ;
      RECT 0.8000 18.2090 104.0460 35.1940 ;
      RECT 0.8000 18.2090 104.0460 35.1940 ;
      RECT 0.8000 18.1650 104.0460 35.1540 ;
      RECT 0.8000 18.1650 104.0460 35.1540 ;
      RECT 0.8000 18.1650 104.0460 35.1540 ;
      RECT 0.0000 9.2950 103.2460 9.2960 ;
      RECT 0.0000 0.8020 103.2460 9.2960 ;
      RECT 0.0000 0.8020 103.2460 9.2960 ;
      RECT 0.0000 0.8020 103.2460 9.2960 ;
      RECT 0.0000 0.8020 104.0460 9.2950 ;
      RECT 0.8000 0.8020 103.2460 16.3030 ;
      RECT 0.8000 0.8020 103.2460 16.3030 ;
      RECT 0.8000 0.8020 103.2460 16.3030 ;
      RECT 84.0600 0.0000 104.0460 9.2950 ;
      RECT 84.0600 0.0000 104.0460 0.8020 ;
      RECT 0.0000 68.7190 104.0460 74.5980 ;
      RECT 0.0000 46.5350 104.0460 52.3970 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.5350 103.2460 53.9600 ;
      RECT 0.8000 46.4960 104.0460 52.3970 ;
      RECT 0.8000 46.4960 104.0460 52.3970 ;
      RECT 0.8000 46.4960 104.0460 52.3970 ;
      RECT 0.8000 46.4960 104.0460 46.5350 ;
      RECT 0.0000 55.3600 104.0460 61.2120 ;
      RECT 0.8000 55.3600 103.2460 65.5020 ;
      RECT 0.8000 55.3600 103.2460 65.5020 ;
      RECT 0.8000 55.3600 103.2460 65.5020 ;
      RECT 0.8000 55.3600 103.2460 65.5020 ;
      RECT 0.8000 55.3600 103.2460 65.5020 ;
      RECT 0.8000 55.3600 103.2460 64.1020 ;
      RECT 0.8000 55.3600 103.2460 64.1020 ;
      RECT 0.8000 55.3600 103.2460 64.1020 ;
      RECT 0.8000 55.3600 103.2460 64.1020 ;
      RECT 0.8000 55.3600 103.2460 64.1020 ;
      RECT 0.8000 55.3600 103.2460 63.7650 ;
      RECT 0.8000 55.3600 103.2460 63.7650 ;
      RECT 0.8000 55.3600 103.2460 63.7650 ;
      RECT 0.8000 55.3600 103.2460 63.7650 ;
      RECT 0.8000 55.3600 103.2460 63.7650 ;
      RECT 0.8000 64.1020 103.2460 74.5980 ;
      RECT 0.8000 64.1020 103.2460 74.5980 ;
      RECT 0.8000 61.2230 103.2460 74.5980 ;
      RECT 0.8000 65.5050 103.2460 68.7190 ;
      RECT 0.8000 64.1020 103.2460 68.7190 ;
      RECT 0.8000 64.1020 103.2460 68.7190 ;
      RECT 0.8000 61.2230 103.2460 68.7190 ;
      RECT 0.8000 65.5050 103.2460 68.7160 ;
      RECT 0.8000 65.5050 103.2460 68.7160 ;
      RECT 0.8000 65.5020 103.2460 68.7160 ;
      RECT 0.8000 65.5020 103.2460 68.7160 ;
      RECT 0.8000 64.1020 103.2460 67.3190 ;
      RECT 0.8000 64.1020 103.2460 67.3190 ;
      RECT 0.8000 61.2230 103.2460 67.3190 ;
      RECT 0.8000 55.3600 103.2460 65.5050 ;
      RECT 0.8000 55.3600 103.2460 65.5050 ;
      RECT 0.8000 55.3600 103.2460 65.5050 ;
      RECT 0.8000 55.3600 103.2460 65.5050 ;
    LAYER PO ;
      RECT 0.0000 0.0000 104.0460 74.5980 ;
    LAYER M3 ;
      RECT 0.0000 68.8190 104.0460 74.5980 ;
      RECT 0.0000 55.4600 104.0460 61.1120 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4230 104.0460 55.4600 ;
      RECT 0.9000 52.3400 103.1460 55.4600 ;
      RECT 0.9000 64.0020 103.1460 74.5980 ;
      RECT 0.9000 64.0020 103.1460 74.5980 ;
      RECT 0.9000 61.1230 103.1460 74.5980 ;
      RECT 0.9000 65.6050 103.1460 68.8190 ;
      RECT 0.9000 64.0020 103.1460 68.8190 ;
      RECT 0.9000 64.0020 103.1460 68.8190 ;
      RECT 0.9000 61.1230 103.1460 68.8190 ;
      RECT 0.9000 65.6050 103.1460 68.8160 ;
      RECT 0.9000 65.6050 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 61.1230 103.1460 67.2190 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 51.7860 0.9000 51.9560 0.9020 ;
      RECT 21.4800 0.0000 22.1680 0.9020 ;
      RECT 0.0000 68.8160 3.0010 68.8190 ;
      RECT 0.0000 65.6020 1.5010 67.2160 ;
      RECT 0.0000 62.7120 0.9000 64.0020 ;
      RECT 51.7860 0.9000 51.9560 1.0510 ;
      RECT 101.0450 61.1120 104.0460 61.1230 ;
      RECT 102.5450 65.6050 104.0460 67.2190 ;
      RECT 103.1460 62.7230 104.0460 63.6650 ;
      RECT 0.0000 52.2970 103.1460 52.3400 ;
      RECT 0.9000 35.0940 103.1460 36.6540 ;
      RECT 0.0000 44.9960 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 104.0460 44.9960 ;
      RECT 0.0000 36.6540 103.1460 36.6940 ;
      RECT 0.0000 46.6350 103.1460 52.3400 ;
      RECT 0.0000 46.6350 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 46.6350 ;
      RECT 0.9000 45.0350 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.0000 16.2030 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 104.0460 16.2030 ;
      RECT 0.0000 0.0000 19.8800 9.1950 ;
      RECT 0.0000 0.0000 19.8800 0.9020 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 10.7960 ;
      RECT 0.9000 9.1960 103.1460 10.7950 ;
      RECT 0.9000 52.3400 103.1460 55.4230 ;
      RECT 0.9000 46.6350 103.1460 55.4230 ;
      RECT 0.0000 18.3090 104.0460 35.0540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 35.0540 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 18.3090 ;
      RECT 0.9000 16.2090 103.1460 18.2650 ;
      RECT 0.0000 9.1950 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 104.0460 9.1950 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 84.1600 0.0000 104.0460 9.1950 ;
      RECT 84.1600 0.0000 104.0460 0.9020 ;
    LAYER M4 ;
      RECT 0.9000 46.6350 103.1460 55.4230 ;
      RECT 0.0000 18.3090 104.0460 35.0540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 35.0540 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 18.3090 ;
      RECT 0.9000 16.2090 103.1460 18.2650 ;
      RECT 0.0000 9.1950 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 104.0460 9.1950 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 84.1600 0.0000 104.0460 9.1950 ;
      RECT 84.1600 0.0000 104.0460 0.9020 ;
      RECT 0.0000 68.8190 104.0460 74.5980 ;
      RECT 0.0000 55.4600 104.0460 61.1120 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 65.6020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4600 103.1460 64.0020 ;
      RECT 0.9000 55.4230 104.0460 55.4600 ;
      RECT 0.9000 52.3400 103.1460 55.4600 ;
      RECT 0.9000 64.0020 103.1460 74.5980 ;
      RECT 0.9000 64.0020 103.1460 74.5980 ;
      RECT 0.9000 61.1230 103.1460 74.5980 ;
      RECT 0.9000 65.6050 103.1460 68.8190 ;
      RECT 0.9000 64.0020 103.1460 68.8190 ;
      RECT 0.9000 64.0020 103.1460 68.8190 ;
      RECT 0.9000 61.1230 103.1460 68.8190 ;
      RECT 0.9000 65.6050 103.1460 68.8160 ;
      RECT 0.9000 65.6050 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 61.1230 103.1460 67.2190 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 0.9000 55.4600 103.1460 65.6050 ;
      RECT 51.7860 0.9000 51.9560 0.9020 ;
      RECT 21.4800 0.0000 22.1680 0.9020 ;
      RECT 0.0000 68.8160 3.0010 68.8190 ;
      RECT 0.0000 65.6020 1.5010 67.2160 ;
      RECT 0.0000 62.7120 0.9000 64.0020 ;
      RECT 51.7860 0.9000 51.9560 1.0510 ;
      RECT 101.0450 61.1120 104.0460 61.1230 ;
      RECT 102.5450 65.6050 104.0460 67.2190 ;
      RECT 103.1460 62.7230 104.0460 63.6650 ;
      RECT 0.0000 52.2970 103.1460 52.3400 ;
      RECT 0.9000 35.0940 103.1460 36.6540 ;
      RECT 0.0000 44.9960 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 104.0460 44.9960 ;
      RECT 0.0000 36.6540 103.1460 36.6940 ;
      RECT 0.0000 46.6350 103.1460 52.3400 ;
      RECT 0.0000 46.6350 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 46.6350 ;
      RECT 0.9000 45.0350 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.0000 16.2030 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 104.0460 16.2030 ;
      RECT 0.0000 0.0000 19.8800 9.1950 ;
      RECT 0.0000 0.0000 19.8800 0.9020 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 10.7960 ;
      RECT 0.9000 9.1960 103.1460 10.7950 ;
      RECT 0.9000 52.3400 103.1460 55.4230 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 104.0460 74.5980 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 104.0460 74.5980 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 104.0460 74.5980 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 104.0460 74.5980 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 104.0460 74.5980 ;
    LAYER M5 ;
      RECT 51.7860 0.9000 51.9560 0.9020 ;
      RECT 0.0000 73.5980 0.7580 74.5980 ;
      RECT 21.4800 0.0000 22.1680 0.9020 ;
      RECT 103.2570 73.5980 104.0460 74.5980 ;
      RECT 0.0000 62.7120 0.9000 64.0020 ;
      RECT 0.0000 65.6020 1.5010 67.2160 ;
      RECT 0.0000 68.8160 3.0010 68.8190 ;
      RECT 0.9000 58.1220 104.0460 61.1230 ;
      RECT 51.7860 0.9000 51.9560 1.0510 ;
      RECT 102.5450 65.6050 104.0460 67.2190 ;
      RECT 103.1460 62.7230 104.0460 63.6650 ;
      RECT 0.0000 16.2030 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 103.1460 16.2090 ;
      RECT 0.0000 10.7960 104.0460 16.2030 ;
      RECT 0.0000 0.0000 19.8800 9.1950 ;
      RECT 0.0000 0.0000 19.8800 0.9020 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 16.2030 ;
      RECT 0.9000 10.7950 104.0460 10.7960 ;
      RECT 0.9000 9.1960 103.1460 10.7950 ;
      RECT 0.9000 18.2650 104.0460 18.3090 ;
      RECT 0.9000 16.2090 103.1460 18.2650 ;
      RECT 0.0000 18.3090 104.0460 35.0540 ;
      RECT 0.9000 35.0940 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 18.3090 103.1460 36.6540 ;
      RECT 0.9000 35.0540 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.3090 104.0460 35.0940 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 18.2650 104.0460 35.0540 ;
      RECT 0.9000 52.3400 103.1460 55.4230 ;
      RECT 0.0000 44.9960 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 103.1460 45.0350 ;
      RECT 0.0000 36.6940 104.0460 44.9960 ;
      RECT 0.0000 36.6540 103.1460 36.6940 ;
      RECT 0.0000 52.2970 103.1460 52.3400 ;
      RECT 0.0000 46.6350 103.1460 52.3400 ;
      RECT 0.0000 46.6350 104.0460 52.2970 ;
      RECT 0.9000 46.6350 103.1460 55.4230 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 52.2970 ;
      RECT 0.9000 46.5960 104.0460 46.6350 ;
      RECT 0.9000 45.0350 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.9000 36.6940 103.1460 46.5960 ;
      RECT 0.0000 9.1950 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 103.1460 9.1960 ;
      RECT 0.0000 0.9020 104.0460 9.1950 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 0.9000 0.9020 103.1460 16.2030 ;
      RECT 84.1600 0.0000 104.0460 9.1950 ;
      RECT 84.1600 0.0000 104.0460 0.9020 ;
      RECT 0.0000 68.8190 104.0460 73.5980 ;
      RECT 0.9000 63.6650 103.1460 64.0020 ;
      RECT 0.0000 55.4600 104.0460 61.1120 ;
      RECT 0.9000 61.1230 103.1460 65.6020 ;
      RECT 0.9000 55.4230 104.0460 55.4600 ;
      RECT 0.9000 52.3400 103.1460 55.4600 ;
      RECT 0.9000 65.6050 103.1460 68.8190 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 65.6020 103.1460 68.8160 ;
      RECT 0.9000 64.0020 103.1460 68.8160 ;
      RECT 0.9000 64.0020 103.1460 68.8160 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
      RECT 0.9000 64.0020 103.1460 67.2190 ;
  END
END SRAMLP2RW32x22

MACRO SRAMLP2RW32x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 132.461 BY 82.535 ;
  SYMMETRY X Y R90 ;

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6320 0.0000 42.8320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6320 0.0000 42.8320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6320 0.0000 42.8320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6320 0.0000 42.8320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6320 0.0000 42.8320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[31]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2640 0.0000 41.4640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2640 0.0000 41.4640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2640 0.0000 41.4640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2640 0.0000 41.4640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2640 0.0000 41.4640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8960 0.0000 40.0960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.8960 0.0000 40.0960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.8960 0.0000 40.0960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.8960 0.0000 40.0960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.8960 0.0000 40.0960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[23]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.5060 0.0020 25.7060 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.5060 0.0020 25.7060 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.5060 0.0020 25.7060 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.5060 0.0020 25.7060 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.5060 0.0020 25.7060 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8480 0.0020 25.0480 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8480 0.0020 25.0480 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8480 0.0020 25.0480 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8480 0.0020 25.0480 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8480 0.0020 25.0480 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.3380 0.0000 81.5380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.3380 0.0000 81.5380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.3380 0.0000 81.5380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.3380 0.0000 81.5380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.3380 0.0000 81.5380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.44356 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.44356 LAYER M4 ;
    ANTENNAMAXAREACAR 15.26851 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 19.40958 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.6880 0.0020 31.8880 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.6880 0.0020 31.8880 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.6880 0.0020 31.8880 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.6880 0.0020 31.8880 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.6880 0.0020 31.8880 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4800 0.0020 23.6800 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4800 0.0020 23.6800 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4800 0.0020 23.6800 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4800 0.0020 23.6800 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4800 0.0020 23.6800 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 1.0572 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 37.92998 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.92998 LAYER M4 ;
    ANTENNAMAXAREACAR 49.12975 LAYER M4 ;
    ANTENNAGATEAREA 1.0572 LAYER M5 ;
    ANTENNAGATEAREA 1.0572 LAYER M6 ;
    ANTENNAGATEAREA 1.0572 LAYER M7 ;
    ANTENNAGATEAREA 1.0572 LAYER M8 ;
    ANTENNAGATEAREA 1.0572 LAYER M9 ;
    ANTENNAGATEAREA 1.0572 LAYER MRDL ;
  END I2[2]

  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.2420 0.0020 28.4420 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.2420 0.0020 28.4420 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.2420 0.0020 28.4420 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.2420 0.0020 28.4420 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.2420 0.0020 28.4420 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[19]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.8750 0.0020 27.0750 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.8750 0.0020 27.0750 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.8750 0.0020 27.0750 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.8750 0.0020 27.0750 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.8750 0.0020 27.0750 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.5840 0.0020 27.7840 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.5840 0.0020 27.7840 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.5840 0.0020 27.7840 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.5840 0.0020 27.7840 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.5840 0.0020 27.7840 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[19]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2160 0.0020 26.4160 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2160 0.0020 26.4160 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2160 0.0020 26.4160 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2160 0.0020 26.4160 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2160 0.0020 26.4160 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.3460 0.0020 32.5460 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.3460 0.0020 32.5460 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.3460 0.0020 32.5460 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.3460 0.0020 32.5460 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.3460 0.0020 32.5460 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.9780 0.0020 31.1780 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.9780 0.0020 31.1780 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.9780 0.0020 31.1780 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.9780 0.0020 31.1780 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.9780 0.0020 31.1780 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.6100 0.0020 29.8100 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.6100 0.0020 29.8100 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.6100 0.0020 29.8100 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.6100 0.0020 29.8100 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.6100 0.0020 29.8100 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[30]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0560 0.0020 33.2560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0560 0.0020 33.2560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0560 0.0020 33.2560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0560 0.0020 33.2560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0560 0.0020 33.2560 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 41.2150 0.2000 41.4150 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 41.2150 0.2000 41.4150 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 41.2150 0.2000 41.4150 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 41.2150 0.2000 41.4150 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 41.2150 0.2000 41.4150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 12.1206 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 10.37596 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.37596 LAYER M3 ;
    ANTENNAMAXAREACAR 27.56834 LAYER M3 ;
    ANTENNAGATEAREA 12.1206 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 11.67182 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.67182 LAYER M4 ;
    ANTENNAMAXAREACAR 673.7904 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A2[4]

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.7700 82.2350 5.0710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.8700 82.2350 4.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.9710 82.2350 3.2710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.0700 82.2350 2.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.1670 82.2350 1.4670 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.6700 82.2350 5.9710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.1700 82.2350 10.4710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.2700 82.2350 9.5710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.3710 82.2350 8.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.4710 82.2350 7.7710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.5710 82.2350 6.8710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.6710 82.2350 14.9710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.7710 82.2350 14.0710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.8700 82.2350 13.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.9710 82.2350 12.2700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.0710 82.2350 11.3710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.5710 82.2350 15.8700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.1700 82.2350 19.4710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.2700 82.2350 18.5710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.3700 82.2350 17.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.4700 82.2350 16.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.8700 82.2350 22.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.9710 82.2350 21.2710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.7700 82.2350 23.0710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.5710 82.2350 24.8700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.6710 82.2350 23.9710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.0710 82.2350 20.3710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.3700 82.2350 26.6700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.2710 82.2350 27.5710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.1700 82.2350 28.4700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.0710 82.2350 29.3710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.4700 82.2350 25.7710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.5710 82.2350 33.8710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.7700 82.2350 32.0710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.9710 82.2350 30.2700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.8710 82.2350 31.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.6700 82.2350 32.9710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.4710 82.2350 34.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.0700 82.2350 38.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.2700 82.2350 36.5710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.1700 82.2350 37.4710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.9700 82.2350 39.2700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.3710 82.2350 35.6700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.4700 82.2350 43.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.8710 82.2350 40.1710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.7700 82.2350 41.0690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.5700 82.2350 42.8700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.6710 82.2350 41.9720 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.9700 82.2350 48.2700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.8710 82.2350 49.1710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.0700 82.2350 47.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.3710 82.2350 44.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.1710 82.2350 46.4720 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.2700 82.2350 45.5690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.4700 82.2350 52.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.7700 82.2350 50.0690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.6710 82.2350 50.9720 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.3710 82.2350 53.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.5700 82.2350 51.8700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.8700 82.2350 58.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.0700 82.2350 56.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.1700 82.2350 55.4700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.2700 82.2350 54.5700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.9710 82.2350 57.2710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.2690 82.2350 63.5690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.3700 82.2350 62.6700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.4700 82.2350 61.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.6700 82.2350 59.9700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.7700 82.2350 59.0700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.5710 82.2350 60.8710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.7690 82.2350 68.0690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.8700 82.2350 67.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.9690 82.2350 66.2690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.0690 82.2350 65.3690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.1700 82.2350 64.4700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.2700 82.2350 72.5700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.3710 82.2350 71.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.4690 82.2350 70.7690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.5690 82.2350 69.8690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.6700 82.2350 68.9700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.7690 82.2350 77.0690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.8700 82.2350 76.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.9700 82.2350 75.2700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.0700 82.2350 74.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.6700 82.2350 77.9700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.1710 82.2350 73.4710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.5690 82.2350 78.8690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.1710 82.2350 82.4710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.2700 82.2350 81.5700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.3710 82.2350 80.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.4690 82.2350 79.7690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.6700 82.2350 86.9700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.5690 82.2350 87.8690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.7690 82.2350 86.0690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.8700 82.2350 85.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.9700 82.2350 84.2700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.0700 82.2350 83.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.3710 82.2350 89.6710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.0700 82.2350 92.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.1700 82.2350 91.4700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.2700 82.2350 90.5700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.4700 82.2350 88.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.5710 82.2350 96.8710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.8700 82.2350 94.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.6700 82.2350 95.9700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.7690 82.2350 95.0690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.9690 82.2350 93.2690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.0700 82.2350 101.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.9690 82.2350 102.2690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.1690 82.2350 100.4690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.2700 82.2350 99.5700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.3700 82.2350 98.6700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.4700 82.2350 97.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.7720 82.2350 104.0720 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.4710 82.2350 106.7710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.5710 82.2350 105.8710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.6710 82.2350 104.9710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.8710 82.2350 103.1710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.9710 82.2350 111.2710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.2710 82.2350 108.5710 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.0700 82.2350 110.3700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.1700 82.2350 109.4700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.3700 82.2350 107.6700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.4700 82.2350 115.7700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.3690 82.2350 116.6690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.5690 82.2350 114.8690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.6700 82.2350 113.9700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.7700 82.2350 113.0700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.8700 82.2350 112.1700 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.1690 82.2350 118.4690 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.8680 82.2350 121.1680 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.9680 82.2350 120.2680 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.0680 82.2350 119.3680 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.2680 82.2350 117.5680 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.3670 82.2350 125.6670 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.6680 82.2350 122.9680 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.4660 82.2350 124.7660 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.5670 82.2350 123.8670 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.2660 82.2350 126.5660 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.1660 82.2350 127.4660 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.0660 82.2350 128.3660 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.9650 82.2350 129.2650 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.7650 82.2350 131.0650 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.8660 82.2350 130.1660 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.7670 82.2350 122.0670 82.5350 ;
    END
  END VSS

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.9200 82.2350 8.2200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.8200 82.2350 9.1190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.7210 82.2350 19.0210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.6210 82.2350 19.9200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.0210 82.2350 124.3210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.9210 82.2350 125.2200 82.5350 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 146.6226 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 146.6226 LAYER M5 ;
  END VDDL

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.451369 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.451369 LAYER M4 ;
    ANTENNAMAXAREACAR 15.48495 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 19.62601 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 3.4200 82.2350 3.7210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.2210 82.2350 5.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.3200 82.2350 4.6200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.5210 82.2350 2.8200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.6200 82.2350 1.9200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.7210 82.2350 10.0200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.0210 82.2350 7.3200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.1210 82.2350 6.4200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.4190 82.2350 12.7200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.5210 82.2350 11.8220 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.6210 82.2350 10.9210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.2200 82.2350 14.5210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.3210 82.2350 13.6200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.8210 82.2350 18.1200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.9210 82.2350 17.2210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.0210 82.2350 16.3210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.1200 82.2350 15.4200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.4210 82.2350 21.7210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.5210 82.2350 20.8210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.1200 82.2350 24.4210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.2210 82.2350 23.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.3200 82.2350 22.6200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.7200 82.2350 28.0210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.6200 82.2350 28.9210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.9200 82.2350 26.2200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.0210 82.2350 25.3210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.8210 82.2350 27.1200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.3210 82.2350 31.6210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.5200 82.2350 29.8210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.1210 82.2350 33.4200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.4200 82.2350 30.7210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.2210 82.2350 32.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.0200 82.2350 34.3210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.7210 82.2350 37.0210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.5210 82.2350 38.8200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.6200 82.2350 37.9200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.9200 82.2350 35.2210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.8210 82.2350 36.1210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.4210 82.2350 39.7220 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.9210 82.2350 44.2220 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.1210 82.2350 42.4210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.0200 82.2350 43.3190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.2200 82.2350 41.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.3200 82.2350 40.6200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.4210 82.2350 48.7220 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.7200 82.2350 46.0200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.6210 82.2350 46.9210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.5200 82.2350 47.8190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.8200 82.2350 45.1200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.9210 82.2350 53.2210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.1210 82.2350 51.4210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.0210 82.2350 52.3200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.3200 82.2350 49.6200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.2200 82.2350 50.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.3200 82.2350 58.6190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.4200 82.2350 57.7190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.6210 82.2350 55.9200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.7200 82.2350 55.0190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.8200 82.2350 54.1190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.5210 82.2350 56.8210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.8200 82.2350 63.1190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.9200 82.2350 62.2190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.0200 82.2350 61.3190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.2210 82.2350 59.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.1210 82.2350 60.4210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.3200 82.2350 67.6190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.4200 82.2350 66.7190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.5190 82.2350 65.8180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.6190 82.2350 64.9180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.7200 82.2350 64.0200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.8210 82.2350 72.1200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.9210 82.2350 71.2200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.0190 82.2350 70.3180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.1190 82.2350 69.4180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.7210 82.2350 73.0210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.2200 82.2350 68.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.3200 82.2350 76.6190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.4200 82.2350 75.7190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.5200 82.2350 74.8190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.6200 82.2350 73.9190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.2200 82.2350 77.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.8210 82.2350 81.1200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.9210 82.2350 80.2200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.0190 82.2350 79.3180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.1190 82.2350 78.4180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.7210 82.2350 82.0210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.1190 82.2350 87.4180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.3200 82.2350 85.6190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.4200 82.2350 84.7190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.5200 82.2350 83.8190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.6200 82.2350 82.9190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.2200 82.2350 86.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.6200 82.2350 91.9190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.7200 82.2350 91.0190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.8200 82.2350 90.1190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.0190 82.2350 88.3180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.9210 82.2350 89.2210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.2190 82.2350 95.5180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.3190 82.2350 94.6180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.5200 82.2350 92.8190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.1210 82.2350 96.4210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.4200 82.2350 93.7200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.5190 82.2350 101.8180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.7200 82.2350 100.0190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.8200 82.2350 99.1190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.9200 82.2350 98.2190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.0200 82.2350 97.3190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.6200 82.2350 100.9200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.0210 82.2350 106.3200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.1210 82.2350 105.4200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.2210 82.2350 104.5200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.4190 82.2350 102.7180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.3220 82.2350 103.6220 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.6200 82.2350 109.9190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.7200 82.2350 109.0190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.9210 82.2350 107.2200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.5210 82.2350 110.8210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.8210 82.2350 108.1210 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.9190 82.2350 116.2180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.1200 82.2350 114.4190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.2200 82.2350 113.5190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.3200 82.2350 112.6190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.4200 82.2350 111.7190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.0200 82.2350 115.3200 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.4180 82.2350 120.7170 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.5180 82.2350 119.8170 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.6180 82.2350 118.9170 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.8190 82.2350 117.1180 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.7190 82.2350 118.0190 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.1170 82.2350 123.4160 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.3180 82.2350 121.6170 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.4160 82.2350 129.7160 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.8160 82.2350 126.1150 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.7160 82.2350 127.0150 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.6160 82.2350 127.9150 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.5160 82.2350 128.8150 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.3150 82.2350 130.6140 82.5350 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.2180 82.2350 122.5180 82.5350 ;
    END
    ANTENNADIFFAREA 10.95167 LAYER M5 ;
    ANTENNADIFFAREA 10.95167 LAYER M6 ;
    ANTENNADIFFAREA 10.95167 LAYER M7 ;
    ANTENNADIFFAREA 10.95167 LAYER M8 ;
    ANTENNADIFFAREA 10.95167 LAYER M9 ;
    ANTENNADIFFAREA 10.95167 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 146.6256 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 146.6256 LAYER M5 ;
  END VDD

  PIN LS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 74.2120 0.2000 74.4120 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 74.2120 0.2000 74.4120 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 74.2120 0.2000 74.4120 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 74.2120 0.2000 74.4120 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 74.2120 0.2000 74.4120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.452025 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.452025 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.944632 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.944632 LAYER M2 ;
    ANTENNAMAXAREACAR 20.93213 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 34.3609 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.40282 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END LS2

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6500 0.0000 93.8500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6500 0.0000 93.8500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6500 0.0000 93.8500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6500 0.0000 93.8500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6500 0.0000 93.8500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 67.2050 132.4610 67.4050 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 67.2050 132.4610 67.4050 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 67.2050 132.4610 67.4050 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 67.2050 132.4610 67.4050 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 67.2050 132.4610 67.4050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2614 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2614 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A1[0]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 50.8990 0.2000 51.0990 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 50.8990 0.2000 51.0990 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 50.8990 0.2000 51.0990 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 50.8990 0.2000 51.0990 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 50.8990 0.2000 51.0990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2773 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2773 LAYER M1 ;
    ANTENNAGATEAREA 10.7373 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 15.25337 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.25337 LAYER M2 ;
    ANTENNAMAXAREACAR 671.9727 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 58.6200 0.2000 58.8200 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 58.6200 0.2000 58.8200 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 58.6200 0.2000 58.8200 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 58.6200 0.2000 58.8200 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 58.6200 0.2000 58.8200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.27676 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27676 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A2[2]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 59.9090 0.2000 60.1090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 59.9090 0.2000 60.1090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 59.9090 0.2000 60.1090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 59.9090 0.2000 60.1090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 59.9090 0.2000 60.1090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.27358 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27358 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A2[1]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 67.2050 0.2000 67.4050 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 67.2050 0.2000 67.4050 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 67.2050 0.2000 67.4050 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 67.2050 0.2000 67.4050 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 67.2050 0.2000 67.4050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.27256 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27256 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A2[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 59.9090 132.4610 60.1090 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 59.9090 132.4610 60.1090 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 59.9090 132.4610 60.1090 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 59.9090 132.4610 60.1090 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 59.9090 132.4610 60.1090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2656 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2656 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A1[1]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.1128 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.72708 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.72708 LAYER M4 ;
    ANTENNAMAXAREACAR 22.91919 LAYER M4 ;
    ANTENNAGATEAREA 67.7022 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 5775.296 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5775.296 LAYER M5 ;
    ANTENNAMAXAREACAR 176.0587 LAYER M5 ;
    ANTENNAGATEAREA 67.7022 LAYER M6 ;
    ANTENNAGATEAREA 67.7022 LAYER M7 ;
    ANTENNAGATEAREA 67.7022 LAYER M8 ;
    ANTENNAGATEAREA 67.7022 LAYER M9 ;
    ANTENNAGATEAREA 67.7022 LAYER MRDL ;
  END CE2

  PIN SD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 70.3100 132.4610 70.5100 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 70.3100 132.4610 70.5100 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 70.3100 132.4610 70.5100 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 70.3100 132.4610 70.5100 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 70.3100 132.4610 70.5100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAGATEAREA 0.2622 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 7.798904 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.798904 LAYER M3 ;
    ANTENNAMAXAREACAR 34.99892 LAYER M3 ;
    ANTENNAGATEAREA 0.2622 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 35.5748 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END SD

  PIN DS2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 71.0040 0.2000 71.2040 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 71.0040 0.2000 71.2040 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 71.0040 0.2000 71.2040 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 71.0040 0.2000 71.2040 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 71.0040 0.2000 71.2040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END DS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.1900 0.0000 21.3900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.1900 0.0000 21.3900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.1900 0.0000 21.3900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.1900 0.0000 21.3900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.1900 0.0000 21.3900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.5178 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.876314 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.876314 LAYER M2 ;
    ANTENNAMAXAREACAR 6.520897 LAYER M2 ;
    ANTENNAGATEAREA 0.5178 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 6.813244 LAYER M3 ;
    ANTENNAGATEAREA 0.5178 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.105571 LAYER M4 ;
    ANTENNAGATEAREA 0.5178 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.39788 LAYER M5 ;
    ANTENNAGATEAREA 0.5178 LAYER M6 ;
    ANTENNAGATEAREA 0.5178 LAYER M7 ;
    ANTENNAGATEAREA 0.5178 LAYER M8 ;
    ANTENNAGATEAREA 0.5178 LAYER M9 ;
    ANTENNAGATEAREA 0.5178 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.2300 0.0000 111.4300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.2300 0.0000 111.4300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.2300 0.0000 111.4300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.2300 0.0000 111.4300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.2300 0.0000 111.4300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.5178 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.882134 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.882134 LAYER M2 ;
    ANTENNAMAXAREACAR 6.532137 LAYER M2 ;
    ANTENNAGATEAREA 0.5178 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 6.824483 LAYER M3 ;
    ANTENNAGATEAREA 0.5178 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.11681 LAYER M4 ;
    ANTENNAGATEAREA 0.5178 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.409118 LAYER M5 ;
    ANTENNAGATEAREA 0.5178 LAYER M6 ;
    ANTENNAGATEAREA 0.5178 LAYER M7 ;
    ANTENNAGATEAREA 0.5178 LAYER M8 ;
    ANTENNAGATEAREA 0.5178 LAYER M9 ;
    ANTENNAGATEAREA 0.5178 LAYER MRDL ;
  END OEB1

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15172 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15172 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.594 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.594 LAYER M2 ;
    ANTENNAMAXAREACAR 11.94867 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.98553 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.02232 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.05904 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 41.2150 132.4610 41.4150 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 41.2150 132.4610 41.4150 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 41.2150 132.4610 41.4150 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 41.2150 132.4610 41.4150 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 41.2150 132.4610 41.4150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M2 ;
    ANTENNAGATEAREA 18.4842 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 16.60857 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.60857 LAYER M3 ;
    ANTENNAMAXAREACAR 16.89077 LAYER M3 ;
    ANTENNAGATEAREA 18.4842 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 27.67812 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.67812 LAYER M4 ;
    ANTENNAMAXAREACAR 1175.378 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A1[4]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0576 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.69846 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.69846 LAYER M4 ;
    ANTENNAMAXAREACAR 42.49996 LAYER M4 ;
    ANTENNAGATEAREA 0.0576 LAYER M5 ;
    ANTENNAGATEAREA 0.0576 LAYER M6 ;
    ANTENNAGATEAREA 0.0576 LAYER M7 ;
    ANTENNAGATEAREA 0.0576 LAYER M8 ;
    ANTENNAGATEAREA 0.0576 LAYER M9 ;
    ANTENNAGATEAREA 0.0576 LAYER MRDL ;
  END CE1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.60414 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.60414 LAYER M2 ;
    ANTENNAMAXAREACAR 12.01807 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 13.05493 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.09171 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.12843 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.8580 0.0000 102.0580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.8580 0.0000 102.0580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.8580 0.0000 102.0580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.8580 0.0000 102.0580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.8580 0.0000 102.0580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.4900 0.0000 100.6900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.4900 0.0000 100.6900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.4900 0.0000 100.6900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.4900 0.0000 100.6900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.4900 0.0000 100.6900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[18]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.1220 0.0000 99.3220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.1220 0.0000 99.3220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.1220 0.0000 99.3220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.1220 0.0000 99.3220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.1220 0.0000 99.3220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.2260 0.0000 103.4260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.2260 0.0000 103.4260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.2260 0.0000 103.4260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.2260 0.0000 103.4260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.2260 0.0000 103.4260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.5940 0.0000 104.7940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.5940 0.0000 104.7940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.5940 0.0000 104.7940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.5940 0.0000 104.7940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.5940 0.0000 104.7940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.5160 0.0020 102.7160 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.5160 0.0020 102.7160 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.5160 0.0020 102.7160 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.5160 0.0020 102.7160 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.5160 0.0020 102.7160 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[17]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.6200 0.0020 106.8200 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.6200 0.0020 106.8200 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.6200 0.0020 106.8200 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.6200 0.0020 106.8200 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.6200 0.0020 106.8200 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.2520 0.0020 105.4520 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.2520 0.0020 105.4520 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.2520 0.0020 105.4520 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.2520 0.0020 105.4520 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.2520 0.0020 105.4520 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[9]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.9620 0.0000 106.1620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.9620 0.0000 106.1620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.9620 0.0000 106.1620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.9620 0.0000 106.1620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.9620 0.0000 106.1620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.3560 0.0020 109.5560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.3560 0.0020 109.5560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.3560 0.0020 109.5560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.3560 0.0020 109.5560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.3560 0.0020 109.5560 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[8]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.7240 0.0020 110.9240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.7240 0.0020 110.9240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.7240 0.0020 110.9240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.7240 0.0020 110.9240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.7240 0.0020 110.9240 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.1340 0.0020 24.3340 0.2020 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.8840 0.0020 104.0840 0.2020 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.9880 0.0020 108.1880 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.1340 0.0020 24.3340 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.9880 0.0020 108.1880 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.1340 0.0020 24.3340 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.9880 0.0020 108.1880 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.1340 0.0020 24.3340 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.1340 0.0020 24.3340 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.6980 0.0000 108.8980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.6980 0.0000 108.8980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.6980 0.0000 108.8980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.6980 0.0000 108.8980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.6980 0.0000 108.8980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.3300 0.0000 107.5300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.3300 0.0000 107.5300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.3300 0.0000 107.5300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.3300 0.0000 107.5300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.3300 0.0000 107.5300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[16]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.0660 0.0000 110.2660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.0660 0.0000 110.2660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.0660 0.0000 110.2660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.0660 0.0000 110.2660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.0660 0.0000 110.2660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN DS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 70.9410 132.4610 71.1410 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 70.9410 132.4610 71.1410 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 70.9410 132.4610 71.1410 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 70.9410 132.4610 71.1410 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 70.9410 132.4610 71.1410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END DS1

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 50.8990 132.4610 51.0990 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 50.8990 132.4610 51.0990 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 50.8990 132.4610 51.0990 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 50.8990 132.4610 51.0990 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 50.8990 132.4610 51.0990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.26614 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26614 LAYER M1 ;
    ANTENNAGATEAREA 17.0643 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 14.09184 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.09184 LAYER M2 ;
    ANTENNAMAXAREACAR 1172.983 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 58.5260 132.4610 58.7260 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 58.5260 132.4610 58.7260 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 58.5260 132.4610 58.7260 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 58.5260 132.4610 58.7260 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 58.5260 132.4610 58.7260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2656 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2656 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END A1[2]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.1480 0.0000 88.3480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.1480 0.0000 88.3480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.1480 0.0000 88.3480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.1480 0.0000 88.3480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.1480 0.0000 88.3480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32655 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32655 LAYER M3 ;
    ANTENNAMAXAREACAR 64.41731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.3640 0.0020 83.5640 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.3640 0.0020 83.5640 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.3640 0.0020 83.5640 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.3640 0.0020 83.5640 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.3640 0.0020 83.5640 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[25]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.5720 0.0020 91.7720 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.5720 0.0020 91.7720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.5720 0.0020 91.7720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.5720 0.0020 91.7720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.5720 0.0020 91.7720 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[29]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.2040 0.0020 90.4040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.2040 0.0020 90.4040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.2040 0.0020 90.4040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.2040 0.0020 90.4040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.2040 0.0020 90.4040 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[22]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.8360 0.0020 89.0360 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.8360 0.0020 89.0360 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.8360 0.0020 89.0360 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.8360 0.0020 89.0360 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.8360 0.0020 89.0360 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[26]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.9140 0.0000 91.1140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.9140 0.0000 91.1140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.9140 0.0000 91.1140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.9140 0.0000 91.1140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.9140 0.0000 91.1140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[29]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.5460 0.0000 89.7460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.5460 0.0000 89.7460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.5460 0.0000 89.7460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.5460 0.0000 89.7460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.5460 0.0000 89.7460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[22]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.3080 0.0020 94.5080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.3080 0.0020 94.5080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.3080 0.0020 94.5080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.3080 0.0020 94.5080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.3080 0.0020 94.5080 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.9400 0.0020 93.1400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.9400 0.0020 93.1400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.9400 0.0020 93.1400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.9400 0.0020 93.1400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.9400 0.0020 93.1400 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[21]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.0180 0.0000 95.2180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.0180 0.0000 95.2180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.0180 0.0000 95.2180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.0180 0.0000 95.2180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.0180 0.0000 95.2180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[27]

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 74.1310 132.4610 74.3310 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 74.1310 132.4610 74.3310 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 74.1310 132.4610 74.3310 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 74.1310 132.4610 74.3310 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 74.1310 132.4610 74.3310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.441885 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.441885 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.959427 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.959427 LAYER M2 ;
    ANTENNAMAXAREACAR 21.22922 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 34.38095 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.42286 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END LS1

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.2820 0.0000 92.4820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.2820 0.0000 92.4820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.2820 0.0000 92.4820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.2820 0.0000 92.4820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.2820 0.0000 92.4820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[21]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.6760 0.0020 95.8760 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.6760 0.0020 95.8760 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.6760 0.0020 95.8760 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.6760 0.0020 95.8760 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.6760 0.0020 95.8760 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[27]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.0440 0.0020 97.2440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.0440 0.0020 97.2440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.0440 0.0020 97.2440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.0440 0.0020 97.2440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.0440 0.0020 97.2440 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[20]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.3860 0.0000 96.5860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.3860 0.0000 96.5860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.3860 0.0000 96.5860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.3860 0.0000 96.5860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.3860 0.0000 96.5860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[20]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.4130 0.0020 98.6130 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.4130 0.0020 98.6130 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.4130 0.0020 98.6130 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.4130 0.0020 98.6130 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.4130 0.0020 98.6130 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[24]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.7540 0.0000 97.9540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.7540 0.0000 97.9540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.7540 0.0000 97.9540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.7540 0.0000 97.9540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.7540 0.0000 97.9540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[24]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.1480 0.0020 101.3480 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.1480 0.0020 101.3480 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.1480 0.0020 101.3480 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.1480 0.0020 101.3480 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.1480 0.0020 101.3480 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[18]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.7800 0.0020 99.9800 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.7800 0.0020 99.9800 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.7800 0.0020 99.9800 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.7800 0.0020 99.9800 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.7800 0.0020 99.9800 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.9880 0.0020 108.1880 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.9880 0.0020 108.1880 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[16]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 103.8840 0.0020 104.0840 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.8840 0.0020 104.0840 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.8840 0.0020 104.0840 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.8840 0.0020 104.0840 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[10]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.4420 0.0000 85.6420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.4420 0.0000 85.6420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.4420 0.0000 85.6420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.4420 0.0000 85.6420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.4420 0.0000 85.6420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.0740 0.0000 84.2740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.0740 0.0000 84.2740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.0740 0.0000 84.2740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.0740 0.0000 84.2740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.0740 0.0000 84.2740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[23]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4680 0.0020 87.6680 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4680 0.0020 87.6680 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4680 0.0020 87.6680 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4680 0.0020 87.6680 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4680 0.0020 87.6680 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[31]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.1000 0.0020 86.3000 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.1000 0.0020 86.3000 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.1000 0.0020 86.3000 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.1000 0.0020 86.3000 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.1000 0.0020 86.3000 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.7320 0.0020 84.9320 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.7320 0.0020 84.9320 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.7320 0.0020 84.9320 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.7320 0.0020 84.9320 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.7320 0.0020 84.9320 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[23]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.0520 0.0020 71.2520 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.0520 0.0020 71.2520 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.0520 0.0020 71.2520 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.0520 0.0020 71.2520 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.0520 0.0020 71.2520 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[14]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.7880 0.0020 73.9880 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.7880 0.0020 73.9880 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.7880 0.0020 73.9880 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.7880 0.0020 73.9880 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.7880 0.0020 73.9880 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[30]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.4200 0.0020 72.6200 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.4200 0.0020 72.6200 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.4200 0.0020 72.6200 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.4200 0.0020 72.6200 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.4200 0.0020 72.6200 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[19]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.4980 0.0000 74.6980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.4980 0.0000 74.6980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.4980 0.0000 74.6980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.4980 0.0000 74.6980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.4980 0.0000 74.6980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.1300 0.0000 73.3300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.1300 0.0000 73.3300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.1300 0.0000 73.3300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.1300 0.0000 73.3300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.1300 0.0000 73.3300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[30]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.7620 0.0000 71.9620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.7620 0.0000 71.9620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.7620 0.0000 71.9620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.7620 0.0000 71.9620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.7620 0.0000 71.9620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[19]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.5240 0.0020 76.7240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.5240 0.0020 76.7240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.5240 0.0020 76.7240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.5240 0.0020 76.7240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.5240 0.0020 76.7240 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.8660 0.0000 76.0660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.8660 0.0000 76.0660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.8660 0.0000 76.0660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.8660 0.0000 76.0660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.8660 0.0000 76.0660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.1560 0.0020 75.3560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.1560 0.0020 75.3560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.1560 0.0020 75.3560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.1560 0.0020 75.3560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.1560 0.0020 75.3560 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.8920 0.0020 78.0920 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.8920 0.0020 78.0920 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.8920 0.0020 78.0920 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.8920 0.0020 78.0920 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.8920 0.0020 78.0920 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.2340 0.0000 77.4340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.2340 0.0000 77.4340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.2340 0.0000 77.4340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.2340 0.0000 77.4340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.2340 0.0000 77.4340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.9960 0.0020 82.1960 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.9960 0.0020 82.1960 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.9960 0.0020 82.1960 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.9960 0.0020 82.1960 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.9960 0.0020 82.1960 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.6280 0.0020 80.8280 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.6280 0.0020 80.8280 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.6280 0.0020 80.8280 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.6280 0.0020 80.8280 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.6280 0.0020 80.8280 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.2600 0.0020 79.4600 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.2600 0.0020 79.4600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.2600 0.0020 79.4600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.2600 0.0020 79.4600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.2600 0.0020 79.4600 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[28]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.3940 0.0000 70.5940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.3940 0.0000 70.5940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.3940 0.0000 70.5940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.3940 0.0000 70.5940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.3940 0.0000 70.5940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.9700 0.0000 80.1700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.9700 0.0000 80.1700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.9700 0.0000 80.1700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.9700 0.0000 80.1700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.9700 0.0000 80.1700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.6020 0.0000 78.8020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.6020 0.0000 78.8020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.6020 0.0000 78.8020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.6020 0.0000 78.8020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.6020 0.0000 78.8020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[28]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.7060 0.0000 82.9060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.7060 0.0000 82.9060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.7060 0.0000 82.9060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.7060 0.0000 82.9060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.7060 0.0000 82.9060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[25]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.8100 0.0000 87.0100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.8100 0.0000 87.0100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.8100 0.0000 87.0100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.8100 0.0000 87.0100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.8100 0.0000 87.0100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[31]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.6800 0.0000 57.8800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.6800 0.0000 57.8800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.6800 0.0000 57.8800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.6800 0.0000 57.8800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.6800 0.0000 57.8800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[17]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.4420 0.0020 62.6420 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.4420 0.0020 62.6420 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.4420 0.0020 62.6420 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.4420 0.0020 62.6420 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.4420 0.0020 62.6420 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.0740 0.0020 61.2740 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.0740 0.0020 61.2740 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.0740 0.0020 61.2740 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.0740 0.0020 61.2740 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.0740 0.0020 61.2740 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.7060 0.0020 59.9060 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.7060 0.0020 59.9060 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.7060 0.0020 59.9060 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.7060 0.0020 59.9060 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.7060 0.0020 59.9060 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.7840 0.0000 61.9840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.7840 0.0000 61.9840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.7840 0.0000 61.9840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.7840 0.0000 61.9840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.7840 0.0000 61.9840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4160 0.0000 60.6160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4160 0.0000 60.6160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4160 0.0000 60.6160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4160 0.0000 60.6160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4160 0.0000 60.6160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0480 0.0000 59.2480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0480 0.0000 59.2480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0480 0.0000 59.2480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0480 0.0000 59.2480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0480 0.0000 59.2480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.3380 0.0020 58.5380 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.3380 0.0020 58.5380 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.3380 0.0020 58.5380 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.3380 0.0020 58.5380 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.3380 0.0020 58.5380 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[17]

  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.8100 0.0020 64.0100 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.8100 0.0020 64.0100 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.8100 0.0020 64.0100 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.8100 0.0020 64.0100 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.8100 0.0020 64.0100 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[16]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1520 0.0000 63.3520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1520 0.0000 63.3520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1520 0.0000 63.3520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1520 0.0000 63.3520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1520 0.0000 63.3520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[16]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.5460 0.0020 66.7460 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.5460 0.0020 66.7460 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.5460 0.0020 66.7460 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.5460 0.0020 66.7460 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.5460 0.0020 66.7460 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.1780 0.0020 65.3780 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.1780 0.0020 65.3780 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.1780 0.0020 65.3780 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.1780 0.0020 65.3780 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.1780 0.0020 65.3780 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.8880 0.0000 66.0880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.8880 0.0000 66.0880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.8880 0.0000 66.0880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.8880 0.0000 66.0880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.8880 0.0000 66.0880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5200 0.0000 64.7200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5200 0.0000 64.7200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5200 0.0000 64.7200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5200 0.0000 64.7200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5200 0.0000 64.7200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.6840 0.0020 69.8840 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.6840 0.0020 69.8840 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.6840 0.0020 69.8840 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.6840 0.0020 69.8840 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.6840 0.0020 69.8840 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.3160 0.0020 68.5160 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.3160 0.0020 68.5160 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.3160 0.0020 68.5160 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.3160 0.0020 68.5160 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.3160 0.0020 68.5160 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.6580 0.0000 67.8580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.6580 0.0000 67.8580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.6580 0.0000 67.8580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.6580 0.0000 67.8580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.6580 0.0000 67.8580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 1.4424 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 44.85651 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 44.85651 LAYER M4 ;
    ANTENNAMAXAREACAR 44.35049 LAYER M4 ;
    ANTENNAGATEAREA 1.4424 LAYER M5 ;
    ANTENNAGATEAREA 1.4424 LAYER M6 ;
    ANTENNAGATEAREA 1.4424 LAYER M7 ;
    ANTENNAGATEAREA 1.4424 LAYER M8 ;
    ANTENNAGATEAREA 1.4424 LAYER M9 ;
    ANTENNAGATEAREA 1.4424 LAYER MRDL ;
  END I1[2]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.0260 0.0000 69.2260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.0260 0.0000 69.2260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.0260 0.0000 69.2260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.0260 0.0000 69.2260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.0260 0.0000 69.2260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.6580 0.0020 44.8580 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.6580 0.0020 44.8580 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.6580 0.0020 44.8580 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.6580 0.0020 44.8580 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.6580 0.0020 44.8580 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[26]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1040 0.0000 48.3040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1040 0.0000 48.3040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1040 0.0000 48.3040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1040 0.0000 48.3040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1040 0.0000 48.3040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3680 0.0000 45.5680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3680 0.0000 45.5680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3680 0.0000 45.5680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3680 0.0000 45.5680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3680 0.0000 45.5680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[22]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7360 0.0000 46.9360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7360 0.0000 46.9360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7360 0.0000 46.9360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7360 0.0000 46.9360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7360 0.0000 46.9360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[29]

  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.7620 0.0020 48.9620 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.7620 0.0020 48.9620 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.7620 0.0020 48.9620 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.7620 0.0020 48.9620 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.7620 0.0020 48.9620 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[21]

  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.3950 0.0020 47.5950 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.3950 0.0020 47.5950 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.3950 0.0020 47.5950 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.3950 0.0020 47.5950 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.3950 0.0020 47.5950 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[29]

  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.0260 0.0020 46.2260 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.0260 0.0020 46.2260 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.0260 0.0020 46.2260 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.0260 0.0020 46.2260 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.0260 0.0020 46.2260 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[22]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.1300 0.0020 50.3300 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.1300 0.0020 50.3300 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.1300 0.0020 50.3300 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.1300 0.0020 50.3300 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.1300 0.0020 50.3300 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[15]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8400 0.0000 51.0400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8400 0.0000 51.0400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8400 0.0000 51.0400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8400 0.0000 51.0400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8400 0.0000 51.0400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[27]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.4720 0.0000 49.6720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.4720 0.0000 49.6720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.4720 0.0000 49.6720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.4720 0.0000 49.6720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.4720 0.0000 49.6720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[15]

  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.8660 0.0020 53.0660 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.8660 0.0020 53.0660 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.8660 0.0020 53.0660 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.8660 0.0020 53.0660 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.8660 0.0020 53.0660 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[20]

  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.4980 0.0020 51.6980 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.4980 0.0020 51.6980 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.4980 0.0020 51.6980 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.4980 0.0020 51.6980 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.4980 0.0020 51.6980 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[27]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.5760 0.0000 53.7760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.5760 0.0000 53.7760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.5760 0.0000 53.7760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.5760 0.0000 53.7760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.5760 0.0000 53.7760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[24]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2080 0.0000 52.4080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2080 0.0000 52.4080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2080 0.0000 52.4080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2080 0.0000 52.4080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2080 0.0000 52.4080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[20]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3120 0.0000 56.5120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3120 0.0000 56.5120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3120 0.0000 56.5120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3120 0.0000 56.5120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3120 0.0000 56.5120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[18]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9440 0.0000 55.1440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9440 0.0000 55.1440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9440 0.0000 55.1440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9440 0.0000 55.1440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9440 0.0000 55.1440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.9700 0.0020 57.1700 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.9700 0.0020 57.1700 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.9700 0.0020 57.1700 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.9700 0.0020 57.1700 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.9700 0.0020 57.1700 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[18]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.6020 0.0020 55.8020 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.6020 0.0020 55.8020 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.6020 0.0020 55.8020 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.6020 0.0020 55.8020 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.6020 0.0020 55.8020 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.2340 0.0020 54.4340 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.2340 0.0020 54.4340 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.2340 0.0020 54.4340 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.2340 0.0020 54.4340 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.2340 0.0020 54.4340 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[24]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3200 0.0020 30.5200 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3200 0.0020 30.5200 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3200 0.0020 30.5200 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3200 0.0020 30.5200 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3200 0.0020 30.5200 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9520 0.0020 29.1520 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9520 0.0020 29.1520 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9520 0.0020 29.1520 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9520 0.0020 29.1520 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9520 0.0020 29.1520 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[30]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.7140 0.0020 33.9140 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.7140 0.0020 33.9140 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.7140 0.0020 33.9140 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.7140 0.0020 33.9140 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.7140 0.0020 33.9140 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.8170 0.0020 38.0170 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.8170 0.0020 38.0170 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.8170 0.0020 38.0170 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.8170 0.0020 38.0170 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.8170 0.0020 38.0170 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4500 0.0020 36.6500 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4500 0.0020 36.6500 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4500 0.0020 36.6500 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4500 0.0020 36.6500 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4500 0.0020 36.6500 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[11]

  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.0820 0.0020 35.2820 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.0820 0.0020 35.2820 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.0820 0.0020 35.2820 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.0820 0.0020 35.2820 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.0820 0.0020 35.2820 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[28]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5280 0.0000 38.7280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5280 0.0000 38.7280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5280 0.0000 38.7280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5280 0.0000 38.7280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5280 0.0000 38.7280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[25]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1600 0.0000 37.3600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1600 0.0000 37.3600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1600 0.0000 37.3600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1600 0.0000 37.3600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1600 0.0000 37.3600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.7920 0.0000 35.9920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.7920 0.0000 35.9920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.7920 0.0000 35.9920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.7920 0.0000 35.9920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.7920 0.0000 35.9920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4240 0.0020 34.6240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4240 0.0020 34.6240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4240 0.0020 34.6240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4240 0.0020 34.6240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4240 0.0020 34.6240 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32124 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32124 LAYER M3 ;
    ANTENNAMAXAREACAR 64.16445 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[28]

  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.2900 0.0020 43.4900 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.2900 0.0020 43.4900 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.2900 0.0020 43.4900 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.2900 0.0020 43.4900 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.2900 0.0020 43.4900 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[31]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.9220 0.0020 42.1220 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.9220 0.0020 42.1220 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.9220 0.0020 42.1220 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.9220 0.0020 42.1220 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.9220 0.0020 42.1220 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5540 0.0020 40.7540 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5540 0.0020 40.7540 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5540 0.0020 40.7540 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5540 0.0020 40.7540 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5540 0.0020 40.7540 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[23]

  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.1860 0.0020 39.3860 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.1860 0.0020 39.3860 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.1860 0.0020 39.3860 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.1860 0.0020 39.3860 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.1860 0.0020 39.3860 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0000 0.0000 44.2000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0000 0.0000 44.2000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0000 0.0000 44.2000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0000 0.0000 44.2000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0000 0.0000 44.2000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.32136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.32136 LAYER M3 ;
    ANTENNAMAXAREACAR 64.17017 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[26]
  OBS
    LAYER M1 ;
      RECT 0.8000 18.1650 132.4610 40.6150 ;
      RECT 0.8000 18.1650 132.4610 40.6150 ;
      RECT 0.8000 18.1650 132.4610 40.6150 ;
      RECT 0.0000 0.0000 20.5900 9.2950 ;
      RECT 0.0000 0.0000 20.5900 9.2950 ;
      RECT 0.0000 0.8000 22.8800 9.2950 ;
      RECT 0.0000 0.8000 22.8800 9.2950 ;
      RECT 0.0000 0.8000 22.8800 0.8020 ;
      RECT 0.0000 10.6960 131.6610 16.3090 ;
      RECT 0.0000 10.6960 131.6610 16.3090 ;
      RECT 0.0000 10.6960 131.6610 16.3090 ;
      RECT 0.0000 10.6960 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 10.6960 ;
      RECT 0.8000 9.2960 131.6610 10.6950 ;
      RECT 0.0000 9.2950 131.6610 9.2960 ;
      RECT 0.0000 0.8020 131.6610 9.2960 ;
      RECT 0.0000 0.8020 131.6610 9.2960 ;
      RECT 0.0000 0.8020 131.6610 9.2960 ;
      RECT 0.0000 0.8020 132.4610 9.2950 ;
      RECT 0.8000 0.8020 131.6610 10.6960 ;
      RECT 0.8000 0.8020 131.6610 10.6960 ;
      RECT 0.8000 0.8020 131.6610 10.6960 ;
      RECT 111.5240 0.8000 132.4610 9.2950 ;
      RECT 111.5240 0.8000 132.4610 9.2950 ;
      RECT 111.5240 0.8000 132.4610 0.8020 ;
      RECT 112.0300 0.0000 132.4610 9.2950 ;
      RECT 112.0300 0.0000 132.4610 9.2950 ;
      RECT 112.0300 0.0000 132.4610 0.8000 ;
      RECT 0.0000 75.0120 132.4610 82.5350 ;
      RECT 0.8000 71.8040 131.6610 82.5350 ;
      RECT 0.8000 71.8040 131.6610 82.5350 ;
      RECT 0.8000 70.4040 131.6610 74.9310 ;
      RECT 0.8000 70.4040 131.6610 74.9310 ;
      RECT 0.8000 70.4040 131.6610 74.9310 ;
      RECT 0.8000 70.4040 131.6610 74.9310 ;
      RECT 0.8000 70.4040 131.6610 74.9310 ;
      RECT 0.8000 70.4040 131.6610 74.9310 ;
      RECT 0.8000 68.0050 131.6610 74.9310 ;
      RECT 0.8000 68.0050 131.6610 74.9310 ;
      RECT 0.8000 68.0050 131.6610 74.9310 ;
      RECT 0.8000 68.0050 131.6610 74.9310 ;
      RECT 0.8000 66.6050 131.6610 74.9310 ;
      RECT 0.8000 66.6050 131.6610 74.9310 ;
      RECT 0.8000 66.6050 131.6610 73.5310 ;
      RECT 0.8000 66.6050 131.6610 73.5310 ;
      RECT 0.8000 66.6050 131.6610 71.8040 ;
      RECT 0.8000 68.0050 131.6610 71.7410 ;
      RECT 0.8000 68.0050 131.6610 71.7410 ;
      RECT 0.8000 68.0050 131.6610 71.7410 ;
      RECT 0.8000 68.0050 131.6610 71.7410 ;
      RECT 0.8000 68.0050 131.6610 71.7410 ;
      RECT 0.8000 68.0050 131.6610 71.7410 ;
      RECT 0.8000 66.6050 131.6610 71.7410 ;
      RECT 0.8000 66.6050 131.6610 71.7410 ;
      RECT 0.8000 66.6050 131.6610 71.7410 ;
      RECT 0.8000 66.6050 131.6610 71.7410 ;
      RECT 67.3460 0.8000 67.7160 0.8020 ;
      RECT 0.0000 68.0050 1.5010 70.4040 ;
      RECT 0.0000 71.8040 1.5010 73.6120 ;
      RECT 21.9900 0.0000 22.8800 0.8000 ;
      RECT 67.3460 0.8000 67.7160 1.1010 ;
      RECT 129.4600 74.9310 132.4610 75.0120 ;
      RECT 130.9600 68.0050 132.4610 69.7100 ;
      RECT 130.9600 71.7410 132.4610 73.5310 ;
      RECT 0.0000 0.0000 20.5900 0.8000 ;
      RECT 0.0000 51.6990 132.4610 57.9260 ;
      RECT 0.0000 60.7090 132.4610 66.6050 ;
      RECT 0.0000 57.9260 131.6610 58.0200 ;
      RECT 0.0000 51.6990 131.6610 58.0200 ;
      RECT 0.0000 51.6990 131.6610 58.0200 ;
      RECT 0.8000 58.0200 131.6610 66.6050 ;
      RECT 0.8000 51.6990 131.6610 66.6050 ;
      RECT 0.8000 58.0200 131.6610 60.7090 ;
      RECT 0.0000 16.3030 131.6610 16.3090 ;
      RECT 0.8000 18.1650 132.4610 18.2430 ;
      RECT 0.8000 16.3090 131.6610 18.1650 ;
      RECT 0.0000 42.0150 132.4610 50.2990 ;
      RECT 0.0000 18.2430 132.4610 40.6150 ;
      RECT 0.8000 50.2990 131.6610 51.6990 ;
      RECT 0.8000 42.0150 131.6610 51.6990 ;
      RECT 0.8000 40.6150 131.6610 50.2990 ;
      RECT 0.8000 40.6150 131.6610 42.0150 ;
    LAYER PO ;
      RECT 0.0000 0.0000 132.4610 82.5350 ;
    LAYER M3 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 71.9040 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 67.4460 0.9000 67.6160 0.9020 ;
      RECT 22.0900 0.0000 22.7800 0.9000 ;
      RECT 0.0000 68.1050 1.5010 70.3040 ;
      RECT 0.0000 71.9040 1.5010 73.5120 ;
      RECT 67.4460 0.9000 67.6160 1.0510 ;
      RECT 129.4600 75.0310 132.4610 75.1120 ;
      RECT 130.9600 68.1050 132.4610 69.6100 ;
      RECT 130.9600 71.8410 132.4610 73.4310 ;
      RECT 0.0000 0.0000 20.4900 0.9000 ;
      RECT 0.0000 51.7990 132.4610 57.8260 ;
      RECT 0.0000 60.8090 132.4610 66.5050 ;
      RECT 0.0000 57.8260 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.9000 57.9200 131.5610 66.5050 ;
      RECT 0.9000 51.7990 131.5610 66.5050 ;
      RECT 0.9000 57.9200 131.5610 60.8090 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 42.1150 132.4610 50.1990 ;
      RECT 0.0000 18.3430 132.4610 40.5150 ;
      RECT 0.9000 50.1990 131.5610 51.7990 ;
      RECT 0.9000 42.1150 131.5610 51.7990 ;
      RECT 0.9000 40.5150 131.5610 50.1990 ;
      RECT 0.9000 40.5150 131.5610 42.1150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 0.9020 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 0.9020 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 0.9000 ;
      RECT 0.0000 75.1120 132.4610 82.5350 ;
      RECT 0.9000 71.9040 131.5610 82.5350 ;
      RECT 0.9000 71.9040 131.5610 82.5350 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
    LAYER M2 ;
      RECT 67.4460 0.9000 67.6160 0.9020 ;
      RECT 0.0000 68.1050 1.5010 70.3040 ;
      RECT 0.0000 71.9040 1.5010 73.5120 ;
      RECT 22.0900 0.0000 22.7800 0.9000 ;
      RECT 67.4460 0.9000 67.6160 1.0510 ;
      RECT 129.4600 75.0310 132.4610 75.1120 ;
      RECT 130.9600 68.1050 132.4610 69.6100 ;
      RECT 130.9600 71.8410 132.4610 73.4310 ;
      RECT 0.0000 0.0000 20.4900 0.9000 ;
      RECT 0.0000 51.7990 132.4610 57.8260 ;
      RECT 0.0000 60.8090 132.4610 66.5050 ;
      RECT 0.0000 57.8260 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.9000 57.9200 131.5610 66.5050 ;
      RECT 0.9000 51.7990 131.5610 66.5050 ;
      RECT 0.9000 57.9200 131.5610 60.8090 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 42.1150 132.4610 50.1990 ;
      RECT 0.0000 18.3430 132.4610 40.5150 ;
      RECT 0.9000 50.1990 131.5610 51.7990 ;
      RECT 0.9000 42.1150 131.5610 51.7990 ;
      RECT 0.9000 40.5150 131.5610 50.1990 ;
      RECT 0.9000 40.5150 131.5610 42.1150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 0.9020 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 0.9020 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 0.9000 ;
      RECT 0.0000 75.1120 132.4610 82.5350 ;
      RECT 0.9000 71.9040 131.5610 82.5350 ;
      RECT 0.9000 71.9040 131.5610 82.5350 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 71.9040 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
    LAYER M4 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 0.9020 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 0.9000 0.9020 131.5610 10.7960 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 0.9020 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 0.9000 ;
      RECT 0.0000 75.1120 132.4610 82.5350 ;
      RECT 0.9000 71.9040 131.5610 82.5350 ;
      RECT 0.9000 71.9040 131.5610 82.5350 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 70.3040 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 71.9040 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 67.4460 0.9000 67.6160 0.9020 ;
      RECT 22.0900 0.0000 22.7800 0.9000 ;
      RECT 0.0000 68.1050 1.5010 70.3040 ;
      RECT 0.0000 71.9040 1.5010 73.5120 ;
      RECT 67.4460 0.9000 67.6160 1.0510 ;
      RECT 129.4600 75.0310 132.4610 75.1120 ;
      RECT 130.9600 68.1050 132.4610 69.6100 ;
      RECT 130.9600 71.8410 132.4610 73.4310 ;
      RECT 0.0000 0.0000 20.4900 0.9000 ;
      RECT 0.0000 51.7990 132.4610 57.8260 ;
      RECT 0.0000 60.8090 132.4610 66.5050 ;
      RECT 0.0000 57.8260 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.9000 57.9200 131.5610 66.5050 ;
      RECT 0.9000 51.7990 131.5610 66.5050 ;
      RECT 0.9000 57.9200 131.5610 60.8090 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 42.1150 132.4610 50.1990 ;
      RECT 0.0000 18.3430 132.4610 40.5150 ;
      RECT 0.9000 50.1990 131.5610 51.7990 ;
      RECT 0.9000 42.1150 131.5610 51.7990 ;
      RECT 0.9000 40.5150 131.5610 50.1990 ;
      RECT 0.9000 40.5150 131.5610 42.1150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 132.4610 82.5350 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 132.4610 82.5350 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 132.4610 82.5350 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 132.4610 82.5350 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 132.4610 82.5350 ;
    LAYER M5 ;
      RECT 67.4460 0.9000 67.6160 0.9020 ;
      RECT 0.0000 81.5350 0.4670 82.5350 ;
      RECT 22.0900 0.0000 22.7800 0.9000 ;
      RECT 131.7650 81.5350 132.4610 82.5350 ;
      RECT 0.0000 71.9040 1.5010 73.5120 ;
      RECT 0.0000 68.1050 1.5010 70.3040 ;
      RECT 67.4460 0.9000 67.6160 1.0510 ;
      RECT 129.4600 75.0310 132.4610 75.1120 ;
      RECT 130.9600 68.1050 132.4610 69.6100 ;
      RECT 130.9600 71.8410 132.4610 73.4310 ;
      RECT 0.0000 0.0000 20.4900 0.9000 ;
      RECT 0.0000 51.7990 132.4610 57.8260 ;
      RECT 0.0000 42.1150 132.4610 50.1990 ;
      RECT 0.9000 50.1990 131.5610 57.8260 ;
      RECT 0.9000 50.1990 131.5610 51.7990 ;
      RECT 0.0000 60.8090 132.4610 66.5050 ;
      RECT 0.0000 57.8260 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.0000 51.7990 131.5610 57.9200 ;
      RECT 0.9000 51.7990 131.5610 66.5050 ;
      RECT 0.9000 57.9200 131.5610 60.8090 ;
      RECT 0.9000 51.7990 131.5610 60.8090 ;
      RECT 0.0000 18.3430 132.4610 40.5150 ;
      RECT 0.9000 40.5150 131.5610 50.1990 ;
      RECT 0.9000 40.5150 131.5610 42.1150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 40.5150 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.0000 20.4900 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 9.1950 ;
      RECT 0.0000 0.9000 22.7800 0.9020 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 0.9000 0.9020 131.5610 16.2030 ;
      RECT 0.9000 0.9020 131.5610 16.2030 ;
      RECT 0.9000 0.9020 131.5610 16.2030 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 9.1950 ;
      RECT 111.6240 0.9000 132.4610 0.9020 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 9.1950 ;
      RECT 112.1300 0.0000 132.4610 0.9000 ;
      RECT 0.0000 75.1120 132.4610 81.5350 ;
      RECT 0.9000 71.9040 131.5610 75.1120 ;
      RECT 0.9000 70.3040 131.5610 75.1120 ;
      RECT 0.9000 68.1050 131.5610 75.0310 ;
      RECT 0.9000 66.5050 131.5610 75.0310 ;
      RECT 0.9000 73.4310 131.5610 73.5120 ;
      RECT 0.9000 70.3040 131.5610 73.5120 ;
      RECT 0.9000 70.3040 131.5610 73.5120 ;
      RECT 0.9000 70.3040 131.5610 73.5120 ;
      RECT 0.9000 68.1050 131.5610 73.5120 ;
      RECT 0.9000 68.1050 131.5610 73.5120 ;
      RECT 0.9000 68.1050 131.5610 73.5120 ;
      RECT 0.9000 68.1050 131.5610 73.5120 ;
      RECT 0.9000 68.1050 131.5610 73.5120 ;
      RECT 0.9000 66.5050 131.5610 73.5120 ;
      RECT 0.9000 66.5050 131.5610 73.5120 ;
      RECT 0.9000 70.3040 131.5610 73.4310 ;
      RECT 0.9000 70.3040 131.5610 73.4310 ;
      RECT 0.9000 68.1050 131.5610 73.4310 ;
      RECT 0.9000 68.1050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 73.4310 ;
      RECT 0.9000 60.8090 131.5610 73.4310 ;
      RECT 0.9000 66.5050 131.5610 71.9040 ;
      RECT 0.9000 60.8090 131.5610 71.9040 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 68.1050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 66.5050 131.5610 71.8410 ;
      RECT 0.9000 60.8090 131.5610 71.8410 ;
  END
END SRAMLP2RW32x32

MACRO SRAMLP2RW32x39
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 150.61 BY 87.143 ;
  SYMMETRY X Y R90 ;

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.1590 0.0000 88.3590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.1590 0.0000 88.3590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.1590 0.0000 88.3590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.1590 0.0000 88.3590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.1590 0.0000 88.3590 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346002 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346002 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.5670 0.0000 87.7670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.5670 0.0000 87.7670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.5670 0.0000 87.7670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.5670 0.0000 87.7670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.5670 0.0000 87.7670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[8]

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 79.6040 0.2000 79.8040 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 79.6040 0.2000 79.8040 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 79.6040 0.2000 79.8040 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 79.6040 0.2000 79.8040 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 79.6040 0.2000 79.8040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 54.5130 150.6100 54.7130 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 54.5130 150.6100 54.7130 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 54.5130 150.6100 54.7130 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 54.5130 150.6100 54.7130 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 54.5130 150.6100 54.7130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 61.8670 150.6100 62.0670 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 61.8670 150.6100 62.0670 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 61.8670 150.6100 62.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 61.8670 150.6100 62.0670 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 61.8670 150.6100 62.0670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 70.8190 150.6100 71.0190 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 70.8190 150.6100 71.0190 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 70.8190 150.6100 71.0190 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 70.8190 150.6100 71.0190 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 70.8190 150.6100 71.0190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.0470 0.0000 110.2470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.0470 0.0000 110.2470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.0470 0.0000 110.2470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.0470 0.0000 110.2470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.0470 0.0000 110.2470 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346002 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346002 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[24]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.4550 0.0000 109.6550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.4550 0.0000 109.6550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.4550 0.0000 109.6550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.4550 0.0000 109.6550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.4550 0.0000 109.6550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[24]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.6780 0.0000 108.8780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.6780 0.0000 108.8780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.6780 0.0000 108.8780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.6780 0.0000 108.8780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.6780 0.0000 108.8780 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343969 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343969 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[23]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.0840 0.0000 108.2840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.0840 0.0000 108.2840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.0840 0.0000 108.2840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.0840 0.0000 108.2840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.0840 0.0000 108.2840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.3130 0.0000 107.5130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.3130 0.0000 107.5130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.3130 0.0000 107.5130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.3130 0.0000 107.5130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.3130 0.0000 107.5130 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.351014 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.351014 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[22]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.7160 0.0000 106.9160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.7160 0.0000 106.9160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.7160 0.0000 106.9160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.7160 0.0000 106.9160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.7160 0.0000 106.9160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.9420 0.0000 106.1420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.9420 0.0000 106.1420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.9420 0.0000 106.1420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.9420 0.0000 106.1420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.9420 0.0000 106.1420 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343484 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343484 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[21]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.3490 0.0000 105.5490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.3490 0.0000 105.5490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.3490 0.0000 105.5490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.3490 0.0000 105.5490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.3490 0.0000 105.5490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.5750 0.0000 104.7750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.5750 0.0000 104.7750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.5750 0.0000 104.7750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.5750 0.0000 104.7750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.5750 0.0000 104.7750 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345947 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345947 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[20]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.9800 0.0000 104.1800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.9800 0.0000 104.1800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.9800 0.0000 104.1800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.9800 0.0000 104.1800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.9800 0.0000 104.1800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[20]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.2060 0.0000 103.4060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.2060 0.0000 103.4060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.2060 0.0000 103.4060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.2060 0.0000 103.4060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.2060 0.0000 103.4060 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[19]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.6160 0.0000 102.8160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.6160 0.0000 102.8160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.6160 0.0000 102.8160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.6160 0.0000 102.8160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.6160 0.0000 102.8160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.8380 0.0000 102.0380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.8380 0.0000 102.0380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.8380 0.0000 102.0380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.8380 0.0000 102.0380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.8380 0.0000 102.0380 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343974 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343974 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[18]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.2430 0.0000 101.4430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.2430 0.0000 101.4430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.2430 0.0000 101.4430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.2430 0.0000 101.4430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.2430 0.0000 101.4430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.4770 0.0000 100.6770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.4770 0.0000 100.6770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.4770 0.0000 100.6770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.4770 0.0000 100.6770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.4770 0.0000 100.6770 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[17]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.1030 0.0000 99.3030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.1030 0.0000 99.3030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.1030 0.0000 99.3030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.1030 0.0000 99.3030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.1030 0.0000 99.3030 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346002 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346002 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[16]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.5110 0.0000 98.7110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.5110 0.0000 98.7110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.5110 0.0000 98.7110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.5110 0.0000 98.7110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.5110 0.0000 98.7110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[16]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.7340 0.0000 97.9340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.7340 0.0000 97.9340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.7340 0.0000 97.9340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.7340 0.0000 97.9340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.7340 0.0000 97.9340 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343969 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343969 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[15]

  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.6440 0.0000 66.8440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.6440 0.0000 66.8440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.6440 0.0000 66.8440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.6440 0.0000 66.8440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.6440 0.0000 66.8440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[32]

  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.8690 0.0000 66.0690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.8690 0.0000 66.0690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.8690 0.0000 66.0690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.8690 0.0000 66.0690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.8690 0.0000 66.0690 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346002 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346002 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[31]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2770 0.0000 65.4770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2770 0.0000 65.4770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2770 0.0000 65.4770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2770 0.0000 65.4770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2770 0.0000 65.4770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[31]

  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5000 0.0000 64.7000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5000 0.0000 64.7000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5000 0.0000 64.7000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5000 0.0000 64.7000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5000 0.0000 64.7000 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343969 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343969 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[30]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.9060 0.0000 64.1060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.9060 0.0000 64.1060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.9060 0.0000 64.1060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.9060 0.0000 64.1060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.9060 0.0000 64.1060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[30]

  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1350 0.0000 63.3350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1350 0.0000 63.3350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1350 0.0000 63.3350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1350 0.0000 63.3350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1350 0.0000 63.3350 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.351014 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.351014 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[29]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.5380 0.0000 62.7380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.5380 0.0000 62.7380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.5380 0.0000 62.7380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.5380 0.0000 62.7380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.5380 0.0000 62.7380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[29]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.1960 0.0000 86.3960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.1960 0.0000 86.3960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.1960 0.0000 86.3960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.1960 0.0000 86.3960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.1960 0.0000 86.3960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.4250 0.0000 85.6250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.4250 0.0000 85.6250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.4250 0.0000 85.6250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.4250 0.0000 85.6250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.4250 0.0000 85.6250 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.351014 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.351014 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[6]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.8280 0.0000 85.0280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.8280 0.0000 85.0280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.8280 0.0000 85.0280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.8280 0.0000 85.0280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.8280 0.0000 85.0280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.0540 0.0000 84.2540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.0540 0.0000 84.2540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.0540 0.0000 84.2540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.0540 0.0000 84.2540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.0540 0.0000 84.2540 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343484 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343484 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[5]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.7370 0.2000 16.9370 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.7370 0.2000 16.9370 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7370 0.2000 16.9370 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.7370 0.2000 16.9370 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.7370 0.2000 16.9370 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.4610 0.0000 83.6610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.4610 0.0000 83.6610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.4610 0.0000 83.6610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.4610 0.0000 83.6610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.4610 0.0000 83.6610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.6870 0.0000 82.8870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.6870 0.0000 82.8870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.6870 0.0000 82.8870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.6870 0.0000 82.8870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.6870 0.0000 82.8870 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345931 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345931 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.0920 0.0000 82.2920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.0920 0.0000 82.2920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.0920 0.0000 82.2920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.0920 0.0000 82.2920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.0920 0.0000 82.2920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[4]

  PIN O2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.4460 0.0000 75.6460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.4460 0.0000 75.6460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.4460 0.0000 75.6460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.4460 0.0000 75.6460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.4460 0.0000 75.6460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[38]

  PIN SD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 75.7020 150.6100 75.9020 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 75.7020 150.6100 75.9020 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 75.7020 150.6100 75.9020 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 75.7020 150.6100 75.9020 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 75.7020 150.6100 75.9020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB2

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 9.7230 150.6100 9.9230 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 9.7230 150.6100 9.9230 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 9.7230 150.6100 9.9230 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 9.7230 150.6100 9.9230 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 9.7230 150.6100 9.9230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB1

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 44.8340 150.6100 45.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 44.8340 150.6100 45.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 44.8340 150.6100 45.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 44.8340 150.6100 45.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 44.8340 150.6100 45.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 44.8320 0.2000 45.0320 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 44.8320 0.2000 45.0320 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 44.8320 0.2000 45.0320 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 44.8320 0.2000 45.0320 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 44.8320 0.2000 45.0320 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[4]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 17.1930 150.6100 17.3930 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 17.1930 150.6100 17.3930 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 17.1930 150.6100 17.3930 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 17.1930 150.6100 17.3930 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 17.1930 150.6100 17.3930 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE1

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.5610 86.8430 7.8610 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.4610 86.8430 8.7600 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.4610 86.8430 17.7610 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.3610 86.8430 18.6600 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.6620 86.8430 141.9620 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.5620 86.8430 142.8610 87.1430 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 129.7710 0.0000 129.9710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.7710 0.0000 129.9710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.7710 0.0000 129.9710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.7710 0.0000 129.9710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 129.7710 0.0000 129.9710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.7900 0.0000 86.9900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.7900 0.0000 86.9900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.7900 0.0000 86.9900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.7900 0.0000 86.9900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.7900 0.0000 86.9900 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343969 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343969 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[7]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 16.7310 150.6100 16.9310 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 16.7310 150.6100 16.9310 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 16.7310 150.6100 16.9310 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 16.7310 150.6100 16.9310 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 16.7310 150.6100 16.9310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 13.8610 86.8430 14.1600 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.2600 86.8430 145.5590 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.7600 86.8430 15.0610 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.1590 86.8430 146.4600 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.9610 86.8430 4.2600 87.1430 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.8600 86.8430 5.1600 87.1430 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 2.6150 86.8420 2.9160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.7150 86.8420 2.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.4160 86.8420 4.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.5160 86.8420 3.8160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.9150 86.8420 9.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.0160 86.8420 8.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.1150 86.8420 7.4150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.2160 86.8420 6.5160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.3150 86.8420 5.6150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.5160 86.8420 12.8160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.4160 86.8420 13.7160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.6150 86.8420 11.9160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.7150 86.8420 11.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.8150 86.8420 10.1160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.8150 86.8420 19.1150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.3150 86.8420 14.6150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.9150 86.8420 18.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.2150 86.8420 15.5160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.0160 86.8420 17.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.1160 86.8420 16.4160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.7160 86.8420 20.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.3150 86.8420 23.6160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.4150 86.8420 22.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.5160 86.8420 21.8160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.6150 86.8420 20.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.2150 86.8420 24.5160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.7150 86.8420 29.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.8150 86.8420 28.1160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.9160 86.8420 27.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.0160 86.8420 26.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.1160 86.8420 25.4160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.5160 86.8420 30.8150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.6160 86.8420 29.9160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.2150 86.8420 33.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.3160 86.8420 32.6160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.4150 86.8420 31.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.7150 86.8420 38.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.8150 86.8420 37.1160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.9150 86.8420 36.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.0150 86.8420 35.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.1160 86.8420 34.4150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.6160 86.8420 38.9160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.4150 86.8420 40.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.5160 86.8420 39.8160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.3150 86.8420 41.6160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.1160 86.8420 43.4150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.2160 86.8420 42.5160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.9150 86.8420 45.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.8160 86.8420 46.1160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.7150 86.8420 47.0150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.6160 86.8420 47.9160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.0150 86.8420 44.3160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.1160 86.8420 52.4160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.3150 86.8420 50.6160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.5160 86.8420 48.8150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.4160 86.8420 49.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.2150 86.8420 51.5160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.0160 86.8420 53.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.6150 86.8420 56.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.8150 86.8420 55.1160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.7150 86.8420 56.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.5150 86.8420 57.8150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.9160 86.8420 54.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.0150 86.8420 62.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.4160 86.8420 58.7160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.3150 86.8420 59.6140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.1150 86.8420 61.4150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.2160 86.8420 60.5170 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.5150 86.8420 66.8150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.4160 86.8420 67.7160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.6150 86.8420 65.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.9160 86.8420 63.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.7160 86.8420 65.0170 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.8150 86.8420 64.1140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.0150 86.8420 71.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.3150 86.8420 68.6140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.2160 86.8420 69.5170 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.9160 86.8420 72.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.1150 86.8420 70.4150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.4150 86.8420 76.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.6150 86.8420 74.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.7150 86.8420 74.0150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.8150 86.8420 73.1150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.5160 86.8420 75.8160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.8140 86.8420 82.1140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.9150 86.8420 81.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.0150 86.8420 80.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.2150 86.8420 78.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.3150 86.8420 77.6150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.1160 86.8420 79.4160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.3140 86.8420 86.6140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.4150 86.8420 85.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.5140 86.8420 84.8140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.6140 86.8420 83.9140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.7150 86.8420 83.0150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.0140 86.8420 89.3140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.1140 86.8420 88.4140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.2150 86.8420 87.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.8150 86.8420 91.1150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.9160 86.8420 90.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.2150 86.8420 96.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.7160 86.8420 92.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.3140 86.8420 95.6140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.4150 86.8420 94.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.5150 86.8420 93.8150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.6150 86.8420 92.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.7160 86.8420 101.0160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.8150 86.8420 100.1150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.9160 86.8420 99.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.0140 86.8420 98.3140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.1140 86.8420 97.4140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.2150 86.8420 105.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.1140 86.8420 106.4140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.3140 86.8420 104.6140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.4150 86.8420 103.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.5150 86.8420 102.8150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.6150 86.8420 101.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.9160 86.8420 108.2160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.6150 86.8420 110.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.7150 86.8420 110.0150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.8150 86.8420 109.1150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.0150 86.8420 107.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.1160 86.8420 115.4160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.4150 86.8420 112.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.2150 86.8420 114.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.3140 86.8420 113.6140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.5140 86.8420 111.8140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.6150 86.8420 119.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.5140 86.8420 120.8140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.7140 86.8420 119.0140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.8150 86.8420 118.1150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.9150 86.8420 117.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.0150 86.8420 116.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.3170 86.8420 122.6170 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.0160 86.8420 125.3160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.1160 86.8420 124.4160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.2160 86.8420 123.5160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.4160 86.8420 121.7160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.5160 86.8420 129.8160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.8160 86.8420 127.1160 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.6150 86.8420 128.9150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.7150 86.8420 128.0150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.9150 86.8420 126.2150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.0150 86.8420 134.3150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.9140 86.8420 135.2140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.1140 86.8420 133.4140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.2150 86.8420 132.5150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.3150 86.8420 131.6150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.4150 86.8420 130.7150 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.7140 86.8420 137.0140 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.4130 86.8420 139.7130 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.5130 86.8420 138.8130 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.6130 86.8420 137.9130 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.8130 86.8420 136.1130 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.9120 86.8420 144.2120 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.2130 86.8420 141.5130 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.0110 86.8420 143.3110 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.1120 86.8420 142.4120 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.8110 86.8420 145.1110 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.7110 86.8420 146.0110 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.6110 86.8420 146.9110 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.5100 86.8420 147.8100 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.3100 86.8420 149.6100 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.4110 86.8420 148.7110 87.1420 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.3120 86.8420 140.6120 87.1420 ;
    END
  END VSS

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 119.0280 0.0000 119.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.0280 0.0000 119.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.0280 0.0000 119.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.0280 0.0000 119.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.0280 0.0000 119.2280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[31]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 119.6220 0.0000 119.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.6220 0.0000 119.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.6220 0.0000 119.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.6220 0.0000 119.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.6220 0.0000 119.8220 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343795 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343795 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[31]

  PIN I1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.3990 0.0000 120.5990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.3990 0.0000 120.5990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.3990 0.0000 120.5990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.3990 0.0000 120.5990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.3990 0.0000 120.5990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[32]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.9910 0.0000 121.1910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.9910 0.0000 121.1910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.9910 0.0000 121.1910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.9910 0.0000 121.1910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.9910 0.0000 121.1910 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346668 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346668 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[32]

  PIN I1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 121.7660 0.0000 121.9660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.7660 0.0000 121.9660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.7660 0.0000 121.9660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 121.7660 0.0000 121.9660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.7660 0.0000 121.9660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[33]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 122.3650 0.0000 122.5650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.3650 0.0000 122.5650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.3650 0.0000 122.5650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 122.3650 0.0000 122.5650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.3650 0.0000 122.5650 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[33]

  PIN I1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 123.1310 0.0000 123.3310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.1310 0.0000 123.3310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.1310 0.0000 123.3310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.1310 0.0000 123.3310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.1310 0.0000 123.3310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[34]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 123.7260 0.0000 123.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.7260 0.0000 123.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.7260 0.0000 123.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.7260 0.0000 123.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.7260 0.0000 123.9260 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343974 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343974 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[34]

  PIN I1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 124.5040 0.0000 124.7040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.5040 0.0000 124.7040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.5040 0.0000 124.7040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 124.5040 0.0000 124.7040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.5040 0.0000 124.7040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[35]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 125.0940 0.0000 125.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.0940 0.0000 125.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.0940 0.0000 125.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 125.0940 0.0000 125.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 125.0940 0.0000 125.2940 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[35]

  PIN I1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 125.8680 0.0000 126.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.8680 0.0000 126.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.8680 0.0000 126.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 125.8680 0.0000 126.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 125.8680 0.0000 126.0680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[36]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 126.4630 0.0000 126.6630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.4630 0.0000 126.6630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.4630 0.0000 126.6630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 126.4630 0.0000 126.6630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 126.4630 0.0000 126.6630 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345931 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345931 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[36]

  PIN I1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 127.2370 0.0000 127.4370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.2370 0.0000 127.4370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.2370 0.0000 127.4370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 127.2370 0.0000 127.4370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 127.2370 0.0000 127.4370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[37]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 127.8300 0.0000 128.0300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.8300 0.0000 128.0300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.8300 0.0000 128.0300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 127.8300 0.0000 128.0300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 127.8300 0.0000 128.0300 0.2000 ;
    END
    ANTENNADIFFAREA 27.27056 LAYER M1 ;
    ANTENNADIFFAREA 27.27056 LAYER M2 ;
    ANTENNADIFFAREA 27.27056 LAYER M3 ;
    ANTENNADIFFAREA 27.27056 LAYER M4 ;
    ANTENNADIFFAREA 27.27056 LAYER M5 ;
    ANTENNADIFFAREA 27.27056 LAYER M6 ;
    ANTENNADIFFAREA 27.27056 LAYER M7 ;
    ANTENNADIFFAREA 27.27056 LAYER M8 ;
    ANTENNADIFFAREA 27.27056 LAYER M9 ;
    ANTENNADIFFAREA 27.27056 LAYER MRDL ;
    ANTENNAGATEAREA 3.9849 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 46.17857 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 46.17857 LAYER M1 ;
    ANTENNAGATEAREA 3.9849 LAYER M2 ;
    ANTENNAGATEAREA 3.9849 LAYER M3 ;
    ANTENNAGATEAREA 3.9849 LAYER M4 ;
    ANTENNAGATEAREA 3.9849 LAYER M5 ;
    ANTENNAGATEAREA 3.9849 LAYER M6 ;
    ANTENNAGATEAREA 3.9849 LAYER M7 ;
    ANTENNAGATEAREA 3.9849 LAYER M8 ;
    ANTENNAGATEAREA 3.9849 LAYER M9 ;
    ANTENNAGATEAREA 3.9849 LAYER MRDL ;
  END O1[37]

  PIN I1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 128.6040 0.0000 128.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.6040 0.0000 128.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.6040 0.0000 128.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 128.6040 0.0000 128.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 128.6040 0.0000 128.8040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[38]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 129.2010 0.0000 129.4010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.2010 0.0000 129.4010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.2010 0.0000 129.4010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.2010 0.0000 129.4010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 129.2010 0.0000 129.4010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O1[38]

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 76.3960 0.2000 76.5960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 76.3960 0.2000 76.5960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 76.3960 0.2000 76.5960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 76.3960 0.2000 76.5960 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 76.3960 0.2000 76.5960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 79.5240 150.6100 79.7240 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 79.5240 150.6100 79.7240 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 79.5240 150.6100 79.7240 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 79.5240 150.6100 79.7240 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 79.5240 150.6100 79.7240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN DS1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 76.3330 150.6100 76.5330 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 76.3330 150.6100 76.5330 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 76.3330 150.6100 76.5330 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 76.3330 150.6100 76.5330 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 76.3330 150.6100 76.5330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS1

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 54.5130 0.2000 54.7130 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 54.5130 0.2000 54.7130 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 54.5130 0.2000 54.7130 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 54.5130 0.2000 54.7130 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 54.5130 0.2000 54.7130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 62.2610 0.2000 62.4610 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 62.2610 0.2000 62.4610 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 62.2610 0.2000 62.4610 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 62.2610 0.2000 62.4610 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 62.2610 0.2000 62.4610 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 63.5230 0.2000 63.7230 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 63.5230 0.2000 63.7230 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 63.5230 0.2000 63.7230 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 63.5230 0.2000 63.7230 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 63.5230 0.2000 63.7230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 70.8190 0.2000 71.0190 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 70.8190 0.2000 71.0190 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 70.8190 0.2000 71.0190 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 70.8190 0.2000 71.0190 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 70.8190 0.2000 71.0190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.4100 63.5230 150.6100 63.7230 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.4100 63.5230 150.6100 63.7230 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.4100 63.5230 150.6100 63.7230 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.4100 63.5230 150.6100 63.7230 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.4100 63.5230 150.6100 63.7230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.2710 0.2000 17.4710 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.2710 0.2000 17.4710 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.2710 0.2000 17.4710 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.2710 0.2000 17.4710 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.2710 0.2000 17.4710 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE2

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.8220 0.0000 111.0220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.8220 0.0000 111.0220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.8220 0.0000 111.0220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.8220 0.0000 111.0220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.8220 0.0000 111.0220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[25]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.4210 0.0000 111.6210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.4210 0.0000 111.6210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.4210 0.0000 111.6210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.4210 0.0000 111.6210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.4210 0.0000 111.6210 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.361727 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.361727 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[25]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 112.1870 0.0000 112.3870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.1870 0.0000 112.3870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.1870 0.0000 112.3870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 112.1870 0.0000 112.3870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.1870 0.0000 112.3870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[26]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 112.7820 0.0000 112.9820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.7820 0.0000 112.9820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.7820 0.0000 112.9820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 112.7820 0.0000 112.9820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.7820 0.0000 112.9820 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343434 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343434 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[26]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 113.5600 0.0000 113.7600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.5600 0.0000 113.7600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.5600 0.0000 113.7600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 113.5600 0.0000 113.7600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.5600 0.0000 113.7600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[27]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 114.1500 0.0000 114.3500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.1500 0.0000 114.3500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.1500 0.0000 114.3500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.1500 0.0000 114.3500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.1500 0.0000 114.3500 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[27]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 114.9240 0.0000 115.1240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.9240 0.0000 115.1240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.9240 0.0000 115.1240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.9240 0.0000 115.1240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.9240 0.0000 115.1240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[28]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 115.5190 0.0000 115.7190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.5190 0.0000 115.7190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.5190 0.0000 115.7190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.5190 0.0000 115.7190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.5190 0.0000 115.7190 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345947 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345947 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[28]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.2930 0.0000 116.4930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.2930 0.0000 116.4930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.2930 0.0000 116.4930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.2930 0.0000 116.4930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.2930 0.0000 116.4930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[29]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.8860 0.0000 117.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.8860 0.0000 117.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.8860 0.0000 117.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.8860 0.0000 117.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.8860 0.0000 117.0860 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343428 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343428 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[29]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 117.6600 0.0000 117.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.6600 0.0000 117.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.6600 0.0000 117.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 117.6600 0.0000 117.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.6600 0.0000 117.8600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[30]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 118.2570 0.0000 118.4570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.2570 0.0000 118.4570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.2570 0.0000 118.4570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 118.2570 0.0000 118.4570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.2570 0.0000 118.4570 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.351014 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.351014 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[30]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.1400 0.0000 97.3400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.1400 0.0000 97.3400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.1400 0.0000 97.3400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.1400 0.0000 97.3400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.1400 0.0000 97.3400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.3690 0.0000 96.5690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.3690 0.0000 96.5690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.3690 0.0000 96.5690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.3690 0.0000 96.5690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.3690 0.0000 96.5690 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.351014 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.351014 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[14]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.7720 0.0000 95.9720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.7720 0.0000 95.9720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.7720 0.0000 95.9720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.7720 0.0000 95.9720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.7720 0.0000 95.9720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.9980 0.0000 95.1980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.9980 0.0000 95.1980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.9980 0.0000 95.1980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.9980 0.0000 95.1980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.9980 0.0000 95.1980 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343484 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343484 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[13]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.4050 0.0000 94.6050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.4050 0.0000 94.6050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.4050 0.0000 94.6050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.4050 0.0000 94.6050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.4050 0.0000 94.6050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6310 0.0000 93.8310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6310 0.0000 93.8310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6310 0.0000 93.8310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6310 0.0000 93.8310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6310 0.0000 93.8310 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345947 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345947 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.0360 0.0000 93.2360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.0360 0.0000 93.2360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.0360 0.0000 93.2360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.0360 0.0000 93.2360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.0360 0.0000 93.2360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[12]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.2620 0.0000 92.4620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.2620 0.0000 92.4620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.2620 0.0000 92.4620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.2620 0.0000 92.4620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.2620 0.0000 92.4620 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[11]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.6720 0.0000 91.8720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.6720 0.0000 91.8720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.6720 0.0000 91.8720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.6720 0.0000 91.8720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.6720 0.0000 91.8720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.8940 0.0000 91.0940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.8940 0.0000 91.0940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.8940 0.0000 91.0940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.8940 0.0000 91.0940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.8940 0.0000 91.0940 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343434 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343434 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[10]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.2990 0.0000 90.4990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.2990 0.0000 90.4990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.2990 0.0000 90.4990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.2990 0.0000 90.4990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.2990 0.0000 90.4990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.5330 0.0000 89.7330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.5330 0.0000 89.7330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.5330 0.0000 89.7330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.5330 0.0000 89.7330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.5330 0.0000 89.7330 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[9]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2340 0.0000 24.4340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2340 0.0000 24.4340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2340 0.0000 24.4340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2340 0.0000 24.4340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2340 0.0000 24.4340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[1]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.7280 0.0000 80.9280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.7280 0.0000 80.9280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.7280 0.0000 80.9280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.7280 0.0000 80.9280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.7280 0.0000 80.9280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[3]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.3180 0.0000 81.5180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.3180 0.0000 81.5180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.3180 0.0000 81.5180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.3180 0.0000 81.5180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.3180 0.0000 81.5180 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[3]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8290 0.0000 25.0290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8290 0.0000 25.0290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8290 0.0000 25.0290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8290 0.0000 25.0290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8290 0.0000 25.0290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[1]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4680 0.0000 23.6680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4680 0.0000 23.6680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4680 0.0000 23.6680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4680 0.0000 23.6680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4680 0.0000 23.6680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[0]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[0]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.1970 0.0000 26.3970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.1970 0.0000 26.3970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.1970 0.0000 26.3970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.1970 0.0000 26.3970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.1970 0.0000 26.3970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[2]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.5660 0.0000 27.7660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.5660 0.0000 27.7660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.5660 0.0000 27.7660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.5660 0.0000 27.7660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.5660 0.0000 27.7660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[3]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9710 0.0000 27.1710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9710 0.0000 27.1710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9710 0.0000 27.1710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9710 0.0000 27.1710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9710 0.0000 27.1710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[3]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6070 0.0000 25.8070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6070 0.0000 25.8070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6070 0.0000 25.8070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6070 0.0000 25.8070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6070 0.0000 25.8070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[2]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5510 0.0000 36.7510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5510 0.0000 36.7510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5510 0.0000 36.7510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5510 0.0000 36.7510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5510 0.0000 36.7510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[10]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.7730 0.0000 35.9730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.7730 0.0000 35.9730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.7730 0.0000 35.9730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.7730 0.0000 35.9730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.7730 0.0000 35.9730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[9]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1780 0.0000 35.3780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1780 0.0000 35.3780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1780 0.0000 35.3780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1780 0.0000 35.3780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1780 0.0000 35.3780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[9]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4120 0.0000 34.6120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4120 0.0000 34.6120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4120 0.0000 34.6120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4120 0.0000 34.6120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4120 0.0000 34.6120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[8]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[8]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0380 0.0000 33.2380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0380 0.0000 33.2380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0380 0.0000 33.2380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0380 0.0000 33.2380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0380 0.0000 33.2380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[7]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4460 0.0000 32.6460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4460 0.0000 32.6460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4460 0.0000 32.6460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4460 0.0000 32.6460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4460 0.0000 32.6460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[7]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.6690 0.0000 31.8690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.6690 0.0000 31.8690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.6690 0.0000 31.8690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.6690 0.0000 31.8690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.6690 0.0000 31.8690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[6]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0750 0.0000 31.2750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0750 0.0000 31.2750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0750 0.0000 31.2750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0750 0.0000 31.2750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0750 0.0000 31.2750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[6]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3040 0.0000 30.5040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3040 0.0000 30.5040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3040 0.0000 30.5040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3040 0.0000 30.5040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3040 0.0000 30.5040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[5]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7070 0.0000 29.9070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7070 0.0000 29.9070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7070 0.0000 29.9070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7070 0.0000 29.9070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7070 0.0000 29.9070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[5]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9330 0.0000 29.1330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9330 0.0000 29.1330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9330 0.0000 29.1330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9330 0.0000 29.1330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9330 0.0000 29.1330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[4]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.2150 0.0000 77.4150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.2150 0.0000 77.4150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.2150 0.0000 77.4150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.2150 0.0000 77.4150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.2150 0.0000 77.4150 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346668 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346668 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[1]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.5890 0.0000 78.7890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.5890 0.0000 78.7890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.5890 0.0000 78.7890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.5890 0.0000 78.7890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.5890 0.0000 78.7890 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[1]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.3550 0.0000 79.5550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.3550 0.0000 79.5550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.3550 0.0000 79.5550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.3550 0.0000 79.5550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.3550 0.0000 79.5550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[2]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.6230 0.0000 76.8230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.6230 0.0000 76.8230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.6230 0.0000 76.8230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.6230 0.0000 76.8230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.6230 0.0000 76.8230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[0]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.9500 0.0000 80.1500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.9500 0.0000 80.1500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.9500 0.0000 80.1500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.9500 0.0000 80.1500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.9500 0.0000 80.1500 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343974 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343974 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O1[2]

  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.4530 0.0000 49.6530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.4530 0.0000 49.6530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.4530 0.0000 49.6530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.4530 0.0000 49.6530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.4530 0.0000 49.6530 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345947 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345947 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[19]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8580 0.0000 49.0580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8580 0.0000 49.0580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8580 0.0000 49.0580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8580 0.0000 49.0580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8580 0.0000 49.0580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[19]

  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.0840 0.0000 48.2840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.0840 0.0000 48.2840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.0840 0.0000 48.2840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.0840 0.0000 48.2840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.0840 0.0000 48.2840 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343454 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343454 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[18]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4940 0.0000 47.6940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4940 0.0000 47.6940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4940 0.0000 47.6940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4940 0.0000 47.6940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4940 0.0000 47.6940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[18]

  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7160 0.0000 46.9160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7160 0.0000 46.9160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7160 0.0000 46.9160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7160 0.0000 46.9160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7160 0.0000 46.9160 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343434 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343434 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[17]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.1210 0.0000 46.3210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.1210 0.0000 46.3210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.1210 0.0000 46.3210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.1210 0.0000 46.3210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.1210 0.0000 46.3210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[17]

  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3550 0.0000 45.5550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3550 0.0000 45.5550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3550 0.0000 45.5550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3550 0.0000 45.5550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3550 0.0000 45.5550 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[16]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[16]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.9820 0.0000 44.1820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.9820 0.0000 44.1820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.9820 0.0000 44.1820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.9820 0.0000 44.1820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.9820 0.0000 44.1820 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34852 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34852 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[15]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3900 0.0000 43.5900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3900 0.0000 43.5900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3900 0.0000 43.5900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3900 0.0000 43.5900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3900 0.0000 43.5900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[15]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6130 0.0000 42.8130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6130 0.0000 42.8130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6130 0.0000 42.8130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6130 0.0000 42.8130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6130 0.0000 42.8130 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34649 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34649 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[14]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0190 0.0000 42.2190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0190 0.0000 42.2190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0190 0.0000 42.2190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0190 0.0000 42.2190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0190 0.0000 42.2190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[14]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2480 0.0000 41.4480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2480 0.0000 41.4480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2480 0.0000 41.4480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2480 0.0000 41.4480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2480 0.0000 41.4480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[13]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6510 0.0000 40.8510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6510 0.0000 40.8510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6510 0.0000 40.8510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6510 0.0000 40.8510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6510 0.0000 40.8510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[13]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8770 0.0000 40.0770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.8770 0.0000 40.0770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.8770 0.0000 40.0770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.8770 0.0000 40.0770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.8770 0.0000 40.0770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[12]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[12]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5100 0.0000 38.7100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5100 0.0000 38.7100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5100 0.0000 38.7100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5100 0.0000 38.7100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5100 0.0000 38.7100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[11]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9150 0.0000 38.1150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9150 0.0000 38.1150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9150 0.0000 38.1150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9150 0.0000 38.1150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9150 0.0000 38.1150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[11]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1410 0.0000 37.3410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1410 0.0000 37.3410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1410 0.0000 37.3410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1410 0.0000 37.3410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1410 0.0000 37.3410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O2[10]

  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.7640 0.0000 61.9640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.7640 0.0000 61.9640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.7640 0.0000 61.9640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.7640 0.0000 61.9640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.7640 0.0000 61.9640 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343484 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343484 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[28]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1710 0.0000 61.3710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1710 0.0000 61.3710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1710 0.0000 61.3710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1710 0.0000 61.3710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1710 0.0000 61.3710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[28]

  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.3970 0.0000 60.5970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.3970 0.0000 60.5970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.3970 0.0000 60.5970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.3970 0.0000 60.5970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.3970 0.0000 60.5970 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345947 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345947 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[27]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.8020 0.0000 60.0020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.8020 0.0000 60.0020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.8020 0.0000 60.0020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.8020 0.0000 60.0020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.8020 0.0000 60.0020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[27]

  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0280 0.0000 59.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0280 0.0000 59.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0280 0.0000 59.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0280 0.0000 59.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0280 0.0000 59.2280 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[26]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.4380 0.0000 58.6380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.4380 0.0000 58.6380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.4380 0.0000 58.6380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.4380 0.0000 58.6380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.4380 0.0000 58.6380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[26]

  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.6600 0.0000 57.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.6600 0.0000 57.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.6600 0.0000 57.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.6600 0.0000 57.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.6600 0.0000 57.8600 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343974 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343974 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[25]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0650 0.0000 57.2650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0650 0.0000 57.2650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0650 0.0000 57.2650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0650 0.0000 57.2650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0650 0.0000 57.2650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[25]

  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.2990 0.0000 56.4990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.2990 0.0000 56.4990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.2990 0.0000 56.4990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.2990 0.0000 56.4990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.2990 0.0000 56.4990 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[24]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[24]

  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9250 0.0000 55.1250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9250 0.0000 55.1250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9250 0.0000 55.1250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9250 0.0000 55.1250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9250 0.0000 55.1250 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.346002 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.346002 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[23]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3330 0.0000 54.5330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.3330 0.0000 54.5330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.3330 0.0000 54.5330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.3330 0.0000 54.5330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.3330 0.0000 54.5330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[23]

  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.5560 0.0000 53.7560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.5560 0.0000 53.7560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.5560 0.0000 53.7560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.5560 0.0000 53.7560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.5560 0.0000 53.7560 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343969 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343969 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[22]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9620 0.0000 53.1620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9620 0.0000 53.1620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9620 0.0000 53.1620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9620 0.0000 53.1620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9620 0.0000 53.1620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[22]

  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.1910 0.0000 52.3910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.1910 0.0000 52.3910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.1910 0.0000 52.3910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.1910 0.0000 52.3910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.1910 0.0000 52.3910 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.351014 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.351014 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[21]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5940 0.0000 51.7940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5940 0.0000 51.7940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5940 0.0000 51.7940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5940 0.0000 51.7940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5940 0.0000 51.7940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[21]

  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8200 0.0000 51.0200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8200 0.0000 51.0200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8200 0.0000 51.0200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8200 0.0000 51.0200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8200 0.0000 51.0200 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343484 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343484 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[20]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.2270 0.0000 50.4270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.2270 0.0000 50.4270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.2270 0.0000 50.4270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.2270 0.0000 50.4270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.2270 0.0000 50.4270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[20]

  PIN I2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.8500 0.0000 75.0500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.8500 0.0000 75.0500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.8500 0.0000 75.0500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.8500 0.0000 75.0500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.8500 0.0000 75.0500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[38]

  PIN O2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.0790 0.0000 74.2790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.0790 0.0000 74.2790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.0790 0.0000 74.2790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.0790 0.0000 74.2790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.0790 0.0000 74.2790 0.2000 ;
    END
    ANTENNADIFFAREA 3.29819 LAYER M1 ;
    ANTENNADIFFAREA 3.29819 LAYER M2 ;
    ANTENNADIFFAREA 3.29819 LAYER M3 ;
    ANTENNADIFFAREA 3.29819 LAYER M4 ;
    ANTENNADIFFAREA 3.29819 LAYER M5 ;
    ANTENNADIFFAREA 3.29819 LAYER M6 ;
    ANTENNADIFFAREA 3.29819 LAYER M7 ;
    ANTENNADIFFAREA 3.29819 LAYER M8 ;
    ANTENNADIFFAREA 3.29819 LAYER M9 ;
    ANTENNADIFFAREA 3.29819 LAYER MRDL ;
    ANTENNAGATEAREA 0.3702 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 7.849064 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 7.849064 LAYER M1 ;
    ANTENNAGATEAREA 0.3702 LAYER M2 ;
    ANTENNAGATEAREA 0.3702 LAYER M3 ;
    ANTENNAGATEAREA 0.3702 LAYER M4 ;
    ANTENNAGATEAREA 0.3702 LAYER M5 ;
    ANTENNAGATEAREA 0.3702 LAYER M6 ;
    ANTENNAGATEAREA 0.3702 LAYER M7 ;
    ANTENNAGATEAREA 0.3702 LAYER M8 ;
    ANTENNAGATEAREA 0.3702 LAYER M9 ;
    ANTENNAGATEAREA 0.3702 LAYER MRDL ;
  END O2[37]

  PIN I2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.4820 0.0000 73.6820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.4820 0.0000 73.6820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.4820 0.0000 73.6820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.4820 0.0000 73.6820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.4820 0.0000 73.6820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[37]

  PIN O2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.7080 0.0000 72.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.7080 0.0000 72.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.7080 0.0000 72.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.7080 0.0000 72.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.7080 0.0000 72.9080 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343484 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343484 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[36]

  PIN I2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.1150 0.0000 72.3150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.1150 0.0000 72.3150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.1150 0.0000 72.3150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.1150 0.0000 72.3150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.1150 0.0000 72.3150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[36]

  PIN O2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.3410 0.0000 71.5410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.3410 0.0000 71.5410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.3410 0.0000 71.5410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.3410 0.0000 71.5410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.3410 0.0000 71.5410 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.345947 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.345947 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[35]

  PIN I2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.7460 0.0000 70.9460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.7460 0.0000 70.9460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.7460 0.0000 70.9460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.7460 0.0000 70.9460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.7460 0.0000 70.9460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[35]

  PIN O2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.9720 0.0000 70.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.9720 0.0000 70.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.9720 0.0000 70.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.9720 0.0000 70.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.9720 0.0000 70.1720 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.34346 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.34346 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[34]

  PIN O2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.6040 0.0000 68.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.6040 0.0000 68.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.6040 0.0000 68.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.6040 0.0000 68.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.6040 0.0000 68.8040 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.343434 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.343434 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[33]

  PIN I2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.3820 0.0000 69.5820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.3820 0.0000 69.5820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.3820 0.0000 69.5820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.3820 0.0000 69.5820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.3820 0.0000 69.5820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[34]

  PIN I2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.0090 0.0000 68.2090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.0090 0.0000 68.2090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.0090 0.0000 68.2090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.0090 0.0000 68.2090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.0090 0.0000 68.2090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[33]

  PIN O2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.2430 0.0000 67.4430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.2430 0.0000 67.4430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.2430 0.0000 67.4430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.2430 0.0000 67.4430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.2430 0.0000 67.4430 0.2000 ;
    END
    ANTENNADIFFAREA 2.176758 LAYER M1 ;
    ANTENNADIFFAREA 2.176758 LAYER M2 ;
    ANTENNADIFFAREA 2.176758 LAYER M3 ;
    ANTENNADIFFAREA 2.176758 LAYER M4 ;
    ANTENNADIFFAREA 2.176758 LAYER M5 ;
    ANTENNADIFFAREA 2.176758 LAYER M6 ;
    ANTENNADIFFAREA 2.176758 LAYER M7 ;
    ANTENNADIFFAREA 2.176758 LAYER M8 ;
    ANTENNADIFFAREA 2.176758 LAYER M9 ;
    ANTENNADIFFAREA 2.176758 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.360887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.360887 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O2[32]
  OBS
    LAYER M2 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 18.1710 ;
      RECT 0.9000 16.0370 149.7100 18.0930 ;
      RECT 0.0000 16.0310 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 150.6100 16.0310 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 10.6240 ;
      RECT 0.9000 9.0240 149.7100 10.6230 ;
      RECT 0.0000 9.0230 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 150.6100 9.0230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 130.6710 0.0000 150.6100 9.0230 ;
      RECT 130.6710 0.0000 150.6100 0.9000 ;
      RECT 0.0000 64.4230 150.6100 70.1190 ;
      RECT 0.0000 55.4130 150.6100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 55.4130 ;
      RECT 0.0000 80.5040 150.6100 87.1430 ;
      RECT 0.9000 77.2960 149.7100 80.4240 ;
      RECT 0.9000 78.8240 149.7100 78.9040 ;
      RECT 0.0000 71.7190 150.6100 75.0020 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 70.1190 149.7100 75.0020 ;
      RECT 0.9000 70.1190 149.7100 71.7190 ;
      RECT 0.9000 62.7670 150.6100 62.8230 ;
      RECT 21.4790 0.0000 22.1690 0.9000 ;
      RECT 0.0000 72.6950 149.7100 75.6960 ;
      RECT 0.0000 77.2960 1.5010 78.9040 ;
      RECT 0.0000 58.5600 149.7100 61.5610 ;
      RECT 149.1090 77.2330 150.6100 78.8240 ;
      RECT 0.9000 80.4240 150.6100 83.4250 ;
      RECT 0.9000 61.5610 149.7100 62.7670 ;
      RECT 0.9000 62.8230 149.7100 65.7680 ;
      RECT 0.0000 45.7320 149.7100 45.7340 ;
      RECT 0.9000 44.1340 149.7100 45.7320 ;
      RECT 0.0000 45.7340 150.6100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 0.0000 19.8790 9.0230 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 18.1710 150.6100 44.1320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 44.1320 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
    LAYER M1 ;
      RECT 0.8000 62.6670 150.6100 62.9230 ;
      RECT 21.3790 0.0000 22.2690 0.8000 ;
      RECT 0.0000 72.7950 149.8100 75.7960 ;
      RECT 0.0000 77.1960 1.5010 79.0040 ;
      RECT 0.0000 58.6600 149.8100 61.6610 ;
      RECT 149.1090 77.1330 150.6100 78.9240 ;
      RECT 0.8000 80.3240 150.6100 83.3250 ;
      RECT 0.8000 61.6610 149.8100 62.6670 ;
      RECT 0.8000 62.9230 149.8100 65.6680 ;
      RECT 0.0000 45.6320 149.8100 45.6340 ;
      RECT 0.8000 44.2340 149.8100 45.6320 ;
      RECT 0.0000 45.6340 150.6100 53.9130 ;
      RECT 0.0000 45.6320 149.8100 53.9130 ;
      RECT 0.0000 45.6320 149.8100 53.9130 ;
      RECT 0.0000 45.6320 149.8100 53.9130 ;
      RECT 0.0000 0.0000 19.9790 9.1230 ;
      RECT 0.0000 0.0000 19.9790 0.8000 ;
      RECT 0.0000 18.0710 150.6100 44.2320 ;
      RECT 0.8000 18.0710 149.8100 45.6320 ;
      RECT 0.8000 18.0710 149.8100 45.6320 ;
      RECT 0.8000 18.0710 149.8100 45.6320 ;
      RECT 0.8000 44.2320 150.6100 44.2340 ;
      RECT 0.8000 18.0710 150.6100 44.2340 ;
      RECT 0.8000 18.0710 150.6100 44.2340 ;
      RECT 0.8000 18.0710 150.6100 44.2340 ;
      RECT 0.8000 17.9930 150.6100 44.2320 ;
      RECT 0.8000 17.9930 150.6100 44.2320 ;
      RECT 0.8000 17.9930 150.6100 44.2320 ;
      RECT 0.8000 17.9930 150.6100 18.0710 ;
      RECT 0.8000 16.1370 149.8100 17.9930 ;
      RECT 0.0000 16.1310 149.8100 16.1370 ;
      RECT 0.0000 10.5240 149.8100 16.1370 ;
      RECT 0.0000 10.5240 149.8100 16.1370 ;
      RECT 0.0000 10.5240 149.8100 16.1370 ;
      RECT 0.0000 10.5240 150.6100 16.1310 ;
      RECT 0.8000 10.5240 149.8100 17.9930 ;
      RECT 0.8000 10.5240 149.8100 17.9930 ;
      RECT 0.8000 10.5240 149.8100 17.9930 ;
      RECT 0.8000 10.5230 150.6100 16.1310 ;
      RECT 0.8000 10.5230 150.6100 16.1310 ;
      RECT 0.8000 10.5230 150.6100 16.1310 ;
      RECT 0.8000 10.5230 150.6100 10.5240 ;
      RECT 0.8000 9.1240 149.8100 10.5230 ;
      RECT 0.0000 9.1230 149.8100 9.1240 ;
      RECT 0.0000 0.8000 149.8100 9.1240 ;
      RECT 0.0000 0.8000 149.8100 9.1240 ;
      RECT 0.0000 0.8000 149.8100 9.1240 ;
      RECT 0.0000 0.8000 150.6100 9.1230 ;
      RECT 0.8000 0.8000 149.8100 10.5230 ;
      RECT 0.8000 0.8000 149.8100 10.5230 ;
      RECT 0.8000 0.8000 149.8100 10.5230 ;
      RECT 130.5710 0.0000 150.6100 9.1230 ;
      RECT 130.5710 0.0000 150.6100 0.8000 ;
      RECT 0.0000 64.3230 150.6100 70.2190 ;
      RECT 0.0000 55.3130 150.6100 61.2670 ;
      RECT 0.8000 53.9130 149.8100 61.2670 ;
      RECT 0.8000 53.9130 149.8100 55.3130 ;
      RECT 0.0000 80.4040 150.6100 87.1430 ;
      RECT 0.8000 77.1960 149.8100 80.3240 ;
      RECT 0.8000 78.9240 149.8100 79.0040 ;
      RECT 0.0000 71.6190 150.6100 75.1020 ;
      RECT 0.8000 77.1330 149.8100 80.3240 ;
      RECT 0.8000 77.1330 149.8100 80.3240 ;
      RECT 0.8000 77.1330 149.8100 80.3240 ;
      RECT 0.8000 77.1330 149.8100 80.3240 ;
      RECT 0.8000 77.1330 149.8100 80.3240 ;
      RECT 0.8000 75.7960 149.8100 80.3240 ;
      RECT 0.8000 75.7960 149.8100 80.3240 ;
      RECT 0.8000 75.7960 149.8100 80.3240 ;
      RECT 0.8000 75.7960 149.8100 80.3240 ;
      RECT 0.8000 75.7960 149.8100 80.3240 ;
      RECT 0.8000 70.2190 149.8100 75.1020 ;
      RECT 0.8000 70.2190 149.8100 71.6190 ;
    LAYER PO ;
      RECT 0.0000 0.0000 150.6100 87.1430 ;
    LAYER M4 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 150.6100 9.0230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 130.6710 0.0000 150.6100 9.0230 ;
      RECT 130.6710 0.0000 150.6100 0.9000 ;
      RECT 0.0000 64.4230 150.6100 70.1190 ;
      RECT 0.0000 55.4130 150.6100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 55.4130 ;
      RECT 0.0000 80.5040 150.6100 87.1430 ;
      RECT 0.9000 77.2960 149.7100 80.4240 ;
      RECT 0.9000 78.8240 149.7100 78.9040 ;
      RECT 0.0000 71.7190 150.6100 75.0020 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 70.1190 149.7100 75.0020 ;
      RECT 0.9000 70.1190 149.7100 71.7190 ;
      RECT 21.4790 0.0000 22.1690 0.9000 ;
      RECT 0.0000 58.5600 149.7100 61.5610 ;
      RECT 0.0000 77.2960 1.5010 78.9040 ;
      RECT 0.0000 72.6950 149.7100 75.6960 ;
      RECT 0.9000 61.5610 149.7100 62.7670 ;
      RECT 0.9000 62.8230 149.7100 65.7680 ;
      RECT 0.9000 62.7670 150.6100 62.8230 ;
      RECT 0.9000 80.4240 150.6100 83.4250 ;
      RECT 149.1090 77.2330 150.6100 78.8240 ;
      RECT 0.0000 45.7320 149.7100 45.7340 ;
      RECT 0.9000 44.1340 149.7100 45.7320 ;
      RECT 0.0000 45.7340 150.6100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 0.0000 19.8790 9.0230 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 18.1710 150.6100 44.1320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 44.1320 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 18.1710 ;
      RECT 0.9000 16.0370 149.7100 18.0930 ;
      RECT 0.0000 16.0310 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 150.6100 16.0310 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 10.6240 ;
      RECT 0.9000 9.0240 149.7100 10.6230 ;
      RECT 0.0000 9.0230 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
    LAYER M3 ;
      RECT 21.4790 0.0000 22.1690 0.9000 ;
      RECT 0.0000 58.5600 149.7100 61.5610 ;
      RECT 0.0000 77.2960 1.5010 78.9040 ;
      RECT 0.0000 72.6950 149.7100 75.6960 ;
      RECT 0.9000 61.5610 149.7100 62.7670 ;
      RECT 0.9000 62.8230 149.7100 65.7680 ;
      RECT 0.9000 62.7670 150.6100 62.8230 ;
      RECT 0.9000 80.4240 150.6100 83.4250 ;
      RECT 149.1090 77.2330 150.6100 78.8240 ;
      RECT 0.0000 45.7320 149.7100 45.7340 ;
      RECT 0.9000 44.1340 149.7100 45.7320 ;
      RECT 0.0000 45.7340 150.6100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 0.0000 19.8790 9.0230 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 18.1710 150.6100 44.1320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 44.1320 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 18.1710 ;
      RECT 0.9000 16.0370 149.7100 18.0930 ;
      RECT 0.0000 16.0310 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 150.6100 16.0310 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 10.6240 ;
      RECT 0.9000 9.0240 149.7100 10.6230 ;
      RECT 0.0000 9.0230 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 150.6100 9.0230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 130.6710 0.0000 150.6100 9.0230 ;
      RECT 130.6710 0.0000 150.6100 0.9000 ;
      RECT 0.0000 64.4230 150.6100 70.1190 ;
      RECT 0.0000 55.4130 150.6100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 55.4130 ;
      RECT 0.0000 80.5040 150.6100 87.1430 ;
      RECT 0.9000 77.2960 149.7100 80.4240 ;
      RECT 0.9000 78.8240 149.7100 78.9040 ;
      RECT 0.0000 71.7190 150.6100 75.0020 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 77.2330 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 70.1190 149.7100 75.0020 ;
      RECT 0.9000 70.1190 149.7100 71.7190 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 150.6100 87.1430 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 150.6100 87.1430 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 150.6100 87.1430 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 150.6100 87.1430 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 150.6100 87.1430 ;
    LAYER M5 ;
      RECT 0.0000 86.1420 1.0150 87.1430 ;
      RECT 21.4790 0.0000 22.1690 0.9000 ;
      RECT 150.3100 86.1420 150.6100 87.1430 ;
      RECT 0.0000 75.0020 3.0010 75.6960 ;
      RECT 0.0000 77.2960 1.5010 78.9040 ;
      RECT 0.0000 58.5600 149.7100 61.5610 ;
      RECT 0.9000 61.5610 149.7100 62.7670 ;
      RECT 0.9000 62.8230 149.7100 65.7680 ;
      RECT 0.9000 62.7670 150.6100 62.8230 ;
      RECT 0.9000 80.4240 150.6100 83.4250 ;
      RECT 149.1090 77.2330 150.6100 78.8240 ;
      RECT 0.0000 0.0000 19.8790 9.0230 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 45.7340 150.6100 53.8130 ;
      RECT 0.9000 9.0240 149.7100 10.6230 ;
      RECT 0.0000 18.1710 150.6100 44.1320 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 53.8130 ;
      RECT 0.0000 45.7320 149.7100 45.7340 ;
      RECT 0.9000 44.1340 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 18.1710 149.7100 45.7320 ;
      RECT 0.9000 44.1320 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.9000 18.1710 150.6100 44.1340 ;
      RECT 0.0000 10.6240 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 16.0310 ;
      RECT 0.9000 10.6230 150.6100 10.6240 ;
      RECT 0.0000 16.0310 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.0000 10.6240 149.7100 16.0370 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 44.1320 ;
      RECT 0.9000 18.0930 150.6100 18.1710 ;
      RECT 0.9000 16.0370 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.9000 10.6240 149.7100 18.0930 ;
      RECT 0.0000 9.0230 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 149.7100 9.0240 ;
      RECT 0.0000 0.9000 150.6100 9.0230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 0.9000 0.9000 149.7100 10.6230 ;
      RECT 130.6710 0.0000 150.6100 9.0230 ;
      RECT 130.6710 0.0000 150.6100 0.9000 ;
      RECT 0.0000 71.7190 150.6100 75.0020 ;
      RECT 0.0000 55.4130 150.6100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 61.1670 ;
      RECT 0.9000 53.8130 149.7100 55.4130 ;
      RECT 0.0000 64.4230 150.6100 70.1190 ;
      RECT 0.9000 64.4230 149.7100 75.0020 ;
      RECT 0.9000 70.1190 149.7100 71.7190 ;
      RECT 0.0000 80.5040 150.6100 86.1420 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 75.6960 149.7100 80.4240 ;
      RECT 0.9000 71.7190 149.7100 78.9040 ;
      RECT 0.9000 71.7190 149.7100 78.9040 ;
      RECT 0.9000 71.7190 149.7100 78.9040 ;
      RECT 0.9000 75.6960 149.7100 78.8240 ;
      RECT 0.9000 75.6960 149.7100 78.8240 ;
      RECT 0.9000 71.7190 149.7100 78.8240 ;
      RECT 0.9000 71.7190 149.7100 78.8240 ;
      RECT 0.9000 71.7190 149.7100 78.8240 ;
      RECT 0.9000 71.7190 149.7100 78.8240 ;
      RECT 0.9000 71.7190 149.7100 78.8240 ;
  END
END SRAMLP2RW32x39

MACRO SRAMLP2RW64x4
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 54.996 BY 90.253 ;
  SYMMETRY X Y R90 ;

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 69.6190 54.9960 69.8190 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 69.6190 54.9960 69.8190 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 69.6190 54.9960 69.8190 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 69.6190 54.9960 69.8190 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 69.6190 54.9960 69.8190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.915408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.915408 LAYER M3 ;
    ANTENNAMAXAREACAR 26.80402 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 30.88966 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 34.97503 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[1]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 76.9180 54.9960 77.1180 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 76.9180 54.9960 77.1180 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 76.9180 54.9960 77.1180 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 76.9180 54.9960 77.1180 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 76.9180 54.9960 77.1180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.915408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.915408 LAYER M3 ;
    ANTENNAMAXAREACAR 26.80402 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 30.88966 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 34.97503 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[0]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 79.0640 54.9960 79.2640 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 79.0640 54.9960 79.2640 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 79.0640 54.9960 79.2640 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 79.0640 54.9960 79.2640 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 79.0640 54.9960 79.2640 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAGATEAREA 0.0792 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 3.274446 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.274446 LAYER M3 ;
    ANTENNAMAXAREACAR 44.36607 LAYER M3 ;
    ANTENNAGATEAREA 0.0792 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 46.252 LAYER M4 ;
    ANTENNAGATEAREA 0.0792 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 48.13779 LAYER M5 ;
    ANTENNAGATEAREA 0.0792 LAYER M6 ;
    ANTENNAGATEAREA 0.0792 LAYER M7 ;
    ANTENNAGATEAREA 0.0792 LAYER M8 ;
    ANTENNAGATEAREA 0.0792 LAYER M9 ;
    ANTENNAGATEAREA 0.0792 LAYER MRDL ;
  END SD

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 79.9100 54.9960 80.1100 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 79.9100 54.9960 80.1100 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 79.9100 54.9960 80.1100 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 79.9100 54.9960 80.1100 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 79.9100 54.9960 80.1100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.241108 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.241108 LAYER M2 ;
    ANTENNAMAXAREACAR 12.76501 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.886454 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.886454 LAYER M3 ;
    ANTENNAMAXAREACAR 64.60874 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 79.34001 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 82.61541 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS1

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 83.0540 54.9960 83.2540 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 83.0540 54.9960 83.2540 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 83.0540 54.9960 83.2540 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 83.0540 54.9960 83.2540 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 83.0540 54.9960 83.2540 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.229765 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.229765 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.938872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.938872 LAYER M2 ;
    ANTENNAMAXAREACAR 20.81647 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 28.17303 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.21535 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.25747 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8540 0.2000 10.0540 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8540 0.2000 10.0540 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8540 0.2000 10.0540 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8540 0.2000 10.0540 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8540 0.2000 10.0540 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.57378 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.57378 LAYER M2 ;
    ANTENNAMAXAREACAR 11.81027 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.84714 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.88394 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.92067 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8680 0.2000 17.0680 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8680 0.2000 17.0680 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8680 0.2000 17.0680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8680 0.2000 17.0680 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8680 0.2000 17.0680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.428089 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.428089 LAYER M4 ;
    ANTENNAMAXAREACAR 13.63436 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.77554 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4290 0.2000 17.6290 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4290 0.2000 17.6290 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4290 0.2000 17.6290 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4290 0.2000 17.6290 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4290 0.2000 17.6290 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.31564 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.31564 LAYER M4 ;
    ANTENNAMAXAREACAR 12.66053 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.09244 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.9660 0.2000 26.1660 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 25.9660 0.2000 26.1660 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9660 0.2000 26.1660 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 25.9660 0.2000 26.1660 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 25.9660 0.2000 26.1660 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.138688 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.138688 LAYER M4 ;
    ANTENNAMAXAREACAR 57.87506 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 65.09029 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[5]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 59.3270 0.2000 59.5270 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 59.3270 0.2000 59.5270 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 59.3270 0.2000 59.5270 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 59.3270 0.2000 59.5270 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 59.3270 0.2000 59.5270 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.917648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.917648 LAYER M3 ;
    ANTENNAMAXAREACAR 26.86522 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.00553 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.14556 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[4]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 60.8520 0.2000 61.0520 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 60.8520 0.2000 61.0520 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 60.8520 0.2000 61.0520 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 60.8520 0.2000 61.0520 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 60.8520 0.2000 61.0520 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.918368 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.918368 LAYER M3 ;
    ANTENNAMAXAREACAR 26.90786 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.04816 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.18819 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 68.1490 0.2000 68.3490 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 68.1490 0.2000 68.3490 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 68.1490 0.2000 68.3490 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 68.1490 0.2000 68.3490 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 68.1490 0.2000 68.3490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.917648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.917648 LAYER M3 ;
    ANTENNAMAXAREACAR 26.86522 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.00553 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.14556 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 76.9670 0.2000 77.1670 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 76.9670 0.2000 77.1670 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 76.9670 0.2000 77.1670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 76.9670 0.2000 77.1670 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 76.9670 0.2000 77.1670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.917648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.917648 LAYER M3 ;
    ANTENNAMAXAREACAR 26.86522 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.00553 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.14556 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 79.8510 0.2000 80.0510 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 79.8510 0.2000 80.0510 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 79.8510 0.2000 80.0510 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 79.8510 0.2000 80.0510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16318 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16318 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.356508 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.356508 LAYER M2 ;
    ANTENNAMAXAREACAR 18.18287 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.110648 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.110648 LAYER M3 ;
    ANTENNAMAXAREACAR 25.79549 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 45.86078 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 49.18232 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS2

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 83.0030 0.2000 83.2030 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 83.0030 0.2000 83.2030 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 83.0030 0.2000 83.2030 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 83.0030 0.2000 83.2030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.328265 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.328265 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.938872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.938872 LAYER M2 ;
    ANTENNAMAXAREACAR 20.81647 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.021 LAYER M3 ;
    ANTENNAMAXAREACAR 28.23019 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.2725 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.31462 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.6860 0.0000 20.8860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.6860 0.0000 20.8860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.6860 0.0000 20.8860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.6860 0.0000 20.8860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.6860 0.0000 20.8860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.081 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56752 LAYER M2 ;
    ANTENNAMAXAREACAR 7.972429 LAYER M2 ;
    ANTENNAGATEAREA 0.081 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 9.843508 LAYER M3 ;
    ANTENNAGATEAREA 0.081 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 11.71446 LAYER M4 ;
    ANTENNAGATEAREA 0.081 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 13.5853 LAYER M5 ;
    ANTENNAGATEAREA 0.081 LAYER M6 ;
    ANTENNAGATEAREA 0.081 LAYER M7 ;
    ANTENNAGATEAREA 0.081 LAYER M8 ;
    ANTENNAGATEAREA 0.081 LAYER M9 ;
    ANTENNAGATEAREA 0.081 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.1180 0.0000 34.3180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.1180 0.0000 34.3180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.1180 0.0000 34.3180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.1180 0.0000 34.3180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.1180 0.0000 34.3180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.081 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.57334 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.57334 LAYER M2 ;
    ANTENNAMAXAREACAR 8.04428 LAYER M2 ;
    ANTENNAGATEAREA 0.081 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 9.915355 LAYER M3 ;
    ANTENNAGATEAREA 0.081 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 11.78631 LAYER M4 ;
    ANTENNAGATEAREA 0.081 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 13.65713 LAYER M5 ;
    ANTENNAGATEAREA 0.081 LAYER M6 ;
    ANTENNAGATEAREA 0.081 LAYER M7 ;
    ANTENNAGATEAREA 0.081 LAYER M8 ;
    ANTENNAGATEAREA 0.081 LAYER M9 ;
    ANTENNAGATEAREA 0.081 LAYER MRDL ;
  END OEB1

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 69.6710 0.2000 69.8710 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 69.6710 0.2000 69.8710 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 69.6710 0.2000 69.8710 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 69.6710 0.2000 69.8710 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 69.6710 0.2000 69.8710 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.9185 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9185 LAYER M3 ;
    ANTENNAMAXAREACAR 26.93643 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.07673 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.21676 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.3850 0.0000 26.5850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.3850 0.0000 26.5850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.3850 0.0000 26.5850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.3850 0.0000 26.5850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.3850 0.0000 26.5850 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.0780 0.0000 27.2780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.0780 0.0000 27.2780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.0780 0.0000 27.2780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.0780 0.0000 27.2780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.0780 0.0000 27.2780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.7530 0.0000 27.9530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.7530 0.0000 27.9530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.7530 0.0000 27.9530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.7530 0.0000 27.9530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.7530 0.0000 27.9530 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.5230 0.0000 29.7230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.5230 0.0000 29.7230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.5230 0.0000 29.7230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.5230 0.0000 29.7230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.5230 0.0000 29.7230 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.8480 0.0010 29.0480 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.8480 0.0010 29.0480 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.8480 0.0010 29.0480 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.8480 0.0010 29.0480 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.8480 0.0010 29.0480 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28572 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28572 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.68795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.9024 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.2160 0.0000 30.4160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.2160 0.0000 30.4160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.2160 0.0000 30.4160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.2160 0.0000 30.4160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.2160 0.0000 30.4160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.8910 0.0000 31.0910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.8910 0.0000 31.0910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.8910 0.0000 31.0910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.8910 0.0000 31.0910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.8910 0.0000 31.0910 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.5840 0.0000 31.7840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.5840 0.0000 31.7840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.5840 0.0000 31.7840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.5840 0.0000 31.7840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.5840 0.0000 31.7840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.2590 0.0000 32.4590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.2590 0.0000 32.4590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.2590 0.0000 32.4590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.2590 0.0000 32.4590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.2590 0.0000 32.4590 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.9520 0.0000 33.1520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.9520 0.0000 33.1520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.9520 0.0000 33.1520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.9520 0.0000 33.1520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.9520 0.0000 33.1520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.6270 0.0000 33.8270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.6270 0.0000 33.8270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.6270 0.0000 33.8270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.6270 0.0000 33.8270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.6270 0.0000 33.8270 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 17.3330 54.9960 17.5330 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 17.3330 54.9960 17.5330 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7950 17.3330 54.9950 17.5330 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7950 17.3330 54.9950 17.5330 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7950 17.3330 54.9950 17.5330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30514 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30514 LAYER M4 ;
    ANTENNAMAXAREACAR 12.70888 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.14079 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 9.8560 54.9960 10.0560 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 9.8560 54.9960 10.0560 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 9.8560 54.9960 10.0560 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 9.8560 54.9960 10.0560 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 9.8560 54.9960 10.0560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.57294 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.57294 LAYER M2 ;
    ANTENNAMAXAREACAR 11.80452 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.84139 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.87819 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.91492 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 16.8630 54.9960 17.0630 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 16.8630 54.9960 17.0630 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 16.8630 54.9960 17.0630 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 16.8630 54.9960 17.0630 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 16.8630 54.9960 17.0630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.428089 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.428089 LAYER M4 ;
    ANTENNAMAXAREACAR 13.63054 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.77172 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 25.9610 54.9960 26.1610 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 25.9610 54.9960 26.1610 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 25.9610 54.9960 26.1610 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 25.9610 54.9960 26.1610 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 25.9610 54.9960 26.1610 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.136551 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.136551 LAYER M4 ;
    ANTENNAMAXAREACAR 57.5985 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 64.81375 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[5]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 59.2810 54.9960 59.4810 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 59.2810 54.9960 59.4810 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 59.2810 54.9960 59.4810 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 59.2810 54.9960 59.4810 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 59.2810 54.9960 59.4810 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.916808 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.916808 LAYER M3 ;
    ANTENNAMAXAREACAR 26.84227 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 30.98258 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.12261 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[4]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 60.8000 54.9960 61.0000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 60.8000 54.9960 61.0000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 60.8000 54.9960 61.0000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 60.8000 54.9960 61.0000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 60.8000 54.9960 61.0000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.916808 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.916808 LAYER M3 ;
    ANTENNAMAXAREACAR 26.84227 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 30.98258 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.12261 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7960 68.0980 54.9960 68.2980 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7960 68.0980 54.9960 68.2980 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7960 68.0980 54.9960 68.2980 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7960 68.0980 54.9960 68.2980 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7960 68.0980 54.9960 68.2980 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.916808 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.916808 LAYER M3 ;
    ANTENNAMAXAREACAR 26.84227 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 30.98258 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.12261 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[2]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.5150 89.9530 6.8150 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.1140 89.9530 19.4140 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.0150 89.9530 20.3150 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.7140 89.9530 50.0140 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.6150 89.9530 50.9150 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.6140 89.9530 5.9150 90.2530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 160.7157 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 160.7157 LAYER M5 ;
  END VDDL

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.0170 0.0000 25.2170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.0170 0.0000 25.2170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.0170 0.0000 25.2170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.0170 0.0000 25.2170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.0170 0.0000 25.2170 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.7100 0.0000 25.9100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.7100 0.0000 25.9100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.7100 0.0000 25.9100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.7100 0.0000 25.9100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.7100 0.0000 25.9100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.3420 0.0000 24.5420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.3420 0.0000 24.5420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.3420 0.0000 24.5420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.3420 0.0000 24.5420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.3420 0.0000 24.5420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.9740 0.0000 23.1740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.9740 0.0000 23.1740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.9740 0.0000 23.1740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.9740 0.0000 23.1740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.9740 0.0000 23.1740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28578 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28578 LAYER M3 ;
    ANTENNAMAXAREACAR 62.47588 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.69081 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.90526 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.6490 0.0000 23.8490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.6490 0.0000 23.8490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.6490 0.0000 23.8490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.6490 0.0000 23.8490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.6490 0.0000 23.8490 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.6150 89.9530 14.9150 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.3140 89.9530 53.6130 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.4150 89.9530 52.7150 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.7150 89.9530 14.0150 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.8140 89.9530 4.1140 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.9150 89.9530 3.2150 90.2530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 160.7151 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 160.7151 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.8640 89.9530 17.1640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.3650 89.9530 48.6650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.9660 89.9530 7.2650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.6640 89.9530 27.9630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.2640 89.9530 49.5630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.1650 89.9530 5.4650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.8640 89.9530 26.1640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.7640 89.9530 27.0640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.0640 89.9530 6.3640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.8650 89.9530 35.1640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.2650 89.9530 13.5640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.9640 89.9530 43.2640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.3640 89.9530 21.6640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.5640 89.9530 46.8640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.9640 89.9530 25.2640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.2650 89.9530 4.5650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.1650 89.9530 50.4660 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.5650 89.9530 28.8660 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.8640 89.9530 8.1650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.3650 89.9530 39.6650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.7650 89.9530 18.0650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.8650 89.9530 44.1650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.2650 89.9530 22.5650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.5640 89.9530 1.8640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.6650 89.9530 45.9660 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.0650 89.9530 24.3660 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.3640 89.9530 3.6650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.7640 89.9530 45.0630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.1640 89.9530 23.4630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.4650 89.9530 2.7640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.2640 89.9530 40.5630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.6640 89.9530 18.9630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.0640 89.9530 42.3640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.4640 89.9530 20.7640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.1650 89.9530 41.4660 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.5620 89.9530 19.8630 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.8650 89.9530 53.1650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.0640 89.9530 51.3640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.2650 89.9530 31.5650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.4640 89.9530 29.7640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.5660 89.9530 10.8660 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.7650 89.9530 9.0650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.7640 89.9530 54.0640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.9640 89.9530 52.2640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.0640 89.9530 33.3640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.1640 89.9530 32.4640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.3640 89.9530 30.6640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.3650 89.9530 12.6650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.4650 89.9530 11.7650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.6650 89.9530 9.9650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.9650 89.9530 34.2640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.5640 89.9530 37.8640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.9640 89.9530 16.2640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.7640 89.9530 36.0650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.1640 89.9530 14.4650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.6640 89.9530 36.9650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.0640 89.9530 15.3650 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.4640 89.9530 38.7640 90.2530 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.4640 89.9530 47.7640 90.2530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 5.49 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1570.698 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1570.698 LAYER M5 ;
    ANTENNAMAXAREACAR 372.4159 LAYER M5 ;
    ANTENNAGATEAREA 5.49 LAYER M6 ;
    ANTENNAGATEAREA 5.49 LAYER M7 ;
    ANTENNAGATEAREA 5.49 LAYER M8 ;
    ANTENNAGATEAREA 5.49 LAYER M9 ;
    ANTENNAGATEAREA 5.49 LAYER MRDL ;
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.8000 16.7330 54.1950 18.1330 ;
      RECT 0.8000 16.2680 54.1960 16.7330 ;
      RECT 0.8000 10.6560 54.1960 16.7330 ;
      RECT 0.8000 10.6560 54.1960 16.7330 ;
      RECT 0.8000 10.6560 54.1960 16.7330 ;
      RECT 0.8000 10.6560 54.1960 16.7330 ;
      RECT 0.0000 0.0000 20.0860 9.2540 ;
      RECT 0.0000 0.0000 20.0860 9.2540 ;
      RECT 0.0000 0.8000 28.2480 9.2540 ;
      RECT 0.0000 0.8000 28.2480 9.2540 ;
      RECT 0.0000 0.8000 28.2480 9.2540 ;
      RECT 0.0000 0.8000 28.2480 0.8010 ;
      RECT 0.8000 9.2560 54.1960 10.6540 ;
      RECT 0.0000 0.8010 54.9960 9.2540 ;
      RECT 0.8000 9.2540 54.9960 9.2560 ;
      RECT 0.8000 0.8010 54.9960 9.2560 ;
      RECT 0.8000 0.8010 54.9960 9.2560 ;
      RECT 0.8000 0.8010 54.9960 9.2560 ;
      RECT 29.6480 0.8000 54.9960 9.2540 ;
      RECT 29.6480 0.8000 54.9960 9.2540 ;
      RECT 29.6480 0.8000 54.9960 9.2540 ;
      RECT 29.6480 0.8000 54.9960 0.8010 ;
      RECT 34.9180 0.0000 54.9960 9.2540 ;
      RECT 34.9180 0.0000 54.9960 9.2540 ;
      RECT 34.9180 0.0000 54.9960 0.8000 ;
      RECT 0.0000 70.4710 54.9960 76.3180 ;
      RECT 0.8000 69.0190 54.1960 69.0710 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 76.3670 54.1960 80.6510 ;
      RECT 0.8000 78.4640 54.1960 79.2510 ;
      RECT 0.8000 80.7100 54.1960 83.8540 ;
      RECT 0.8000 80.6510 54.1960 83.8540 ;
      RECT 0.8000 80.6510 54.1960 83.8540 ;
      RECT 0.8000 79.2510 54.1960 83.8540 ;
      RECT 0.8000 79.2510 54.1960 83.8540 ;
      RECT 0.8000 76.3670 54.1960 83.8540 ;
      RECT 0.8000 76.3670 54.1960 83.8540 ;
      RECT 0.8000 80.6510 54.1960 83.8030 ;
      RECT 0.8000 80.6510 54.1960 83.8030 ;
      RECT 0.8000 80.6510 54.1960 83.8030 ;
      RECT 0.8000 80.6510 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 83.8030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.8000 76.3670 54.1960 82.4030 ;
      RECT 0.0000 61.6520 54.9960 67.4980 ;
      RECT 0.0000 26.7660 54.9960 58.6810 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.7270 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 58.6810 54.1960 67.4980 ;
      RECT 0.8000 60.0810 54.1960 60.1270 ;
      RECT 0.8000 26.7610 54.9960 58.6810 ;
      RECT 0.8000 26.7610 54.9960 58.6810 ;
      RECT 0.8000 26.7610 54.9960 58.6810 ;
      RECT 0.8000 26.7610 54.9960 26.7660 ;
      RECT 53.4950 80.7100 54.9960 82.4540 ;
      RECT 0.0000 80.6510 1.5010 82.4030 ;
      RECT 0.0000 77.7670 0.8000 79.2510 ;
      RECT 54.1960 77.7180 54.9960 78.4640 ;
      RECT 0.0000 73.4200 54.1960 76.3670 ;
      RECT 0.0000 73.3660 54.9960 73.4200 ;
      RECT 0.8000 70.4190 54.9960 73.3660 ;
      RECT 0.8000 69.0710 54.1960 70.4190 ;
      RECT 0.0000 69.0190 54.1960 69.0710 ;
      RECT 0.0000 68.9490 54.9960 69.0190 ;
      RECT 0.8000 68.8980 54.9960 68.9490 ;
      RECT 0.8000 67.5490 54.1960 68.8980 ;
      RECT 0.0000 64.5480 54.1960 67.5490 ;
      RECT 51.9950 61.6000 54.9960 61.6520 ;
      RECT 0.0000 60.1270 0.8000 60.2520 ;
      RECT 54.1960 60.0810 54.9960 60.2000 ;
      RECT 0.0000 58.6810 3.0010 58.7270 ;
      RECT 21.4860 0.0000 22.3740 0.8000 ;
      RECT 0.0000 0.0000 20.0860 0.8000 ;
      RECT 0.0000 83.8540 54.9960 90.2530 ;
      RECT 0.0000 83.8030 54.1960 83.8540 ;
      RECT 0.0000 25.3610 54.1960 25.3660 ;
      RECT 0.0000 18.2290 54.1960 25.3660 ;
      RECT 0.0000 18.2290 54.1960 25.3660 ;
      RECT 0.0000 18.2290 54.1960 25.3660 ;
      RECT 0.0000 18.2290 54.9960 25.3610 ;
      RECT 0.8000 25.3660 54.1960 26.7610 ;
      RECT 0.8000 18.2290 54.1960 26.7610 ;
      RECT 0.8000 18.2290 54.1960 26.7610 ;
      RECT 0.8000 18.2290 54.1960 26.7610 ;
      RECT 0.8000 18.1330 54.9960 25.3610 ;
      RECT 0.8000 18.1330 54.9960 25.3610 ;
      RECT 0.8000 18.1330 54.9960 25.3610 ;
      RECT 0.8000 18.1330 54.9960 25.3610 ;
      RECT 0.8000 18.1330 54.9960 18.2290 ;
      RECT 0.0000 16.2630 54.1960 16.2680 ;
      RECT 0.0000 10.6560 54.1960 16.2680 ;
      RECT 0.0000 10.6560 54.1960 16.2680 ;
      RECT 0.0000 10.6560 54.1960 16.2680 ;
      RECT 0.0000 10.6560 54.1960 16.2680 ;
      RECT 0.0000 10.6560 54.9960 16.2630 ;
      RECT 0.0000 10.6540 54.1960 16.2630 ;
      RECT 0.0000 10.6540 54.1960 16.2630 ;
      RECT 0.0000 10.6540 54.1960 16.2630 ;
      RECT 0.0000 10.6540 54.1960 10.6560 ;
      RECT 0.8000 10.6560 54.1950 25.3610 ;
      RECT 0.8000 10.6560 54.1950 25.3610 ;
      RECT 0.8000 10.6560 54.1950 25.3610 ;
      RECT 0.8000 10.6560 54.1950 25.3610 ;
    LAYER PO ;
      RECT 0.0000 0.0000 54.9960 90.2530 ;
    LAYER M2 ;
      RECT 0.9000 16.1680 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.0000 25.2610 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.9960 25.2610 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 26.8660 ;
      RECT 0.9000 25.2660 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 18.2330 54.9960 18.3290 ;
      RECT 0.0000 0.9010 54.9960 9.1540 ;
      RECT 0.9000 9.1540 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 0.9010 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 0.9000 ;
      RECT 0.9000 79.1510 54.0960 90.2530 ;
      RECT 0.9000 79.1510 54.0960 90.2530 ;
      RECT 0.9000 80.8100 54.0960 83.9540 ;
      RECT 0.9000 79.1510 54.0960 83.9540 ;
      RECT 0.9000 79.1510 54.0960 83.9540 ;
      RECT 0.9000 80.8100 54.0960 83.9030 ;
      RECT 0.9000 80.8100 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 82.3030 54.0960 82.3540 ;
      RECT 0.9000 79.1510 54.0960 82.3540 ;
      RECT 0.9000 79.1510 54.0960 82.3540 ;
      RECT 0.9000 80.8100 54.0960 82.3030 ;
      RECT 0.0000 70.5710 54.9960 76.2180 ;
      RECT 0.9000 70.5190 54.9960 70.5710 ;
      RECT 0.9000 67.4490 54.0960 70.5710 ;
      RECT 0.9000 76.2670 54.0960 90.2530 ;
      RECT 0.9000 76.2670 54.0960 90.2530 ;
      RECT 0.9000 76.2670 54.0960 83.9540 ;
      RECT 0.9000 76.2670 54.0960 82.3540 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 78.3640 54.0960 79.1510 ;
      RECT 21.5860 0.0000 22.2740 0.9000 ;
      RECT 53.4950 80.8100 54.9960 82.3540 ;
      RECT 0.0000 73.2660 54.0960 76.2670 ;
      RECT 0.0000 80.7510 1.5010 82.3030 ;
      RECT 54.0960 77.8180 54.9960 78.3640 ;
      RECT 0.0000 77.8670 0.9000 79.1510 ;
      RECT 0.0000 0.0000 19.9860 0.9000 ;
      RECT 0.0000 61.7520 54.9960 67.3980 ;
      RECT 0.0000 26.8660 54.9960 58.5810 ;
      RECT 0.0000 58.5810 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.0960 58.6270 ;
      RECT 0.9000 61.7000 54.9960 67.3980 ;
      RECT 0.9000 58.6270 54.0960 67.3980 ;
      RECT 0.9000 61.7000 54.9960 61.7520 ;
      RECT 0.9000 58.6270 54.0960 61.7000 ;
      RECT 0.9000 26.8660 54.0960 61.7000 ;
      RECT 0.0000 67.3980 54.0960 67.4490 ;
      RECT 0.0000 61.7520 54.0960 67.4490 ;
      RECT 0.9000 67.4490 54.0960 70.5190 ;
      RECT 0.9000 61.7520 54.0960 70.5190 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 0.9010 ;
      RECT 0.9000 9.1560 54.0960 10.7540 ;
      RECT 0.0000 83.9540 54.9960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 83.9540 ;
      RECT 0.9000 82.3540 54.0960 83.9030 ;
      RECT 0.0000 16.1630 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.9960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 10.7560 ;
      RECT 0.9000 16.6330 54.0950 18.2330 ;
    LAYER M3 ;
      RECT 53.4950 80.8100 54.9960 82.3540 ;
      RECT 0.0000 83.9540 54.9960 90.2530 ;
      RECT 0.0000 0.0000 19.9860 0.9000 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 0.9010 ;
      RECT 0.9000 9.1560 54.0960 10.7540 ;
      RECT 0.0000 16.1630 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.9960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 10.7560 ;
      RECT 0.9000 16.6330 54.0950 18.2330 ;
      RECT 0.9000 16.1680 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.9000 10.7560 54.0960 16.6330 ;
      RECT 0.0000 67.3980 54.0960 67.4490 ;
      RECT 0.0000 61.7520 54.0960 67.4490 ;
      RECT 0.0000 61.7520 54.9960 67.3980 ;
      RECT 0.9000 67.4490 54.0960 70.5190 ;
      RECT 0.9000 61.7520 54.0960 70.5190 ;
      RECT 0.0000 25.2610 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.9960 25.2610 ;
      RECT 0.9000 25.2660 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 10.7560 54.0950 25.2610 ;
      RECT 0.9000 18.2330 54.9960 18.3290 ;
      RECT 0.0000 58.5810 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.9960 58.5810 ;
      RECT 0.9000 61.7000 54.9960 67.3980 ;
      RECT 0.9000 58.6270 54.0960 67.3980 ;
      RECT 0.9000 61.7000 54.9960 61.7520 ;
      RECT 0.9000 58.6270 54.0960 61.7000 ;
      RECT 0.9000 26.8660 54.0960 61.7000 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 26.8660 ;
      RECT 0.0000 0.9010 54.9960 9.1540 ;
      RECT 0.9000 9.1540 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 0.9010 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 0.9000 ;
      RECT 0.0000 70.5710 54.9960 76.2180 ;
      RECT 0.9000 70.5190 54.9960 76.2180 ;
      RECT 0.9000 67.4490 54.0960 76.2180 ;
      RECT 0.9000 70.5190 54.9960 70.5710 ;
      RECT 0.0000 78.3640 54.0960 83.9540 ;
      RECT 0.0000 77.8670 54.0960 82.3540 ;
      RECT 0.0000 78.3640 54.0960 82.3540 ;
      RECT 0.0000 77.8670 54.0960 82.3540 ;
      RECT 0.0000 77.8670 54.0960 82.3540 ;
      RECT 21.5860 0.0000 22.2740 0.9000 ;
      RECT 0.0000 73.2660 54.0960 76.2670 ;
      RECT 0.9000 77.8180 54.9960 78.3640 ;
      RECT 0.9000 78.3640 54.0960 79.2680 ;
      RECT 0.9000 76.2670 54.0960 77.8180 ;
    LAYER M5 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 78.3640 54.0960 79.1510 ;
      RECT 54.7640 89.2530 54.9960 90.2530 ;
      RECT 0.0000 89.2530 0.8640 90.2530 ;
      RECT 21.5860 0.0000 22.2740 0.9000 ;
      RECT 21.5860 0.0000 22.2740 0.9010 ;
      RECT 0.0000 77.8670 0.9000 79.1510 ;
      RECT 0.0000 80.7510 1.5010 82.3030 ;
      RECT 0.0000 73.2660 54.0960 76.2670 ;
      RECT 53.4950 80.8100 54.9960 82.3540 ;
      RECT 54.0960 77.8180 54.9960 78.3640 ;
      RECT 0.0000 0.0000 19.9860 0.9000 ;
      RECT 0.0000 67.3980 54.0960 67.4490 ;
      RECT 0.9000 67.4490 54.0960 70.5190 ;
      RECT 0.0000 61.7520 54.0960 67.4490 ;
      RECT 0.0000 61.7520 54.9960 67.3980 ;
      RECT 0.9000 61.7520 54.0960 70.5190 ;
      RECT 0.9000 61.7000 54.9960 67.3980 ;
      RECT 0.9000 58.6270 54.0960 67.3980 ;
      RECT 0.9000 61.7000 54.9960 61.7520 ;
      RECT 0.9000 58.6270 54.0960 61.7000 ;
      RECT 0.0000 83.9540 54.9960 89.2530 ;
      RECT 0.0000 83.9030 54.0960 83.9540 ;
      RECT 0.9000 82.3540 54.0960 83.9030 ;
      RECT 0.0000 58.5810 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.9960 58.5810 ;
      RECT 0.9000 26.8660 54.0960 61.7000 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 26.8660 ;
      RECT 0.9000 25.2660 54.0960 26.8610 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.9000 28.1480 0.9010 ;
      RECT 0.9000 9.1560 54.0960 10.7540 ;
      RECT 0.0000 25.2610 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.9960 25.2610 ;
      RECT 0.0000 16.1630 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.9960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 10.7560 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 10.7560 54.0960 25.2610 ;
      RECT 0.9000 10.7560 54.0960 25.2610 ;
      RECT 0.9000 10.7560 54.0960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 18.3290 ;
      RECT 0.9000 16.1680 54.0960 18.2330 ;
      RECT 0.0000 0.9010 54.9960 9.1540 ;
      RECT 0.9000 9.1540 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 0.9010 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 0.9000 ;
      RECT 0.9000 80.8100 54.0960 83.9540 ;
      RECT 0.9000 80.7510 54.0960 83.9540 ;
      RECT 0.9000 80.7510 54.0960 83.9540 ;
      RECT 0.9000 79.1510 54.0960 83.9540 ;
      RECT 0.9000 79.1510 54.0960 83.9540 ;
      RECT 0.9000 80.8100 54.0960 83.9030 ;
      RECT 0.9000 80.8100 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 82.3030 54.0960 82.3540 ;
      RECT 0.0000 70.5710 54.9960 76.2180 ;
      RECT 0.9000 70.5190 54.9960 70.5710 ;
      RECT 0.9000 67.4490 54.0960 70.5710 ;
      RECT 0.9000 76.2670 54.0960 83.9540 ;
      RECT 0.9000 76.2670 54.0960 83.9540 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 83.9030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
    LAYER M4 ;
      RECT 21.5860 0.0000 22.2740 0.9010 ;
      RECT 21.5860 0.0000 22.2740 0.9000 ;
      RECT 0.0000 77.8670 0.9000 79.1510 ;
      RECT 0.0000 80.7510 1.5010 82.3030 ;
      RECT 0.0000 73.2660 54.0960 76.2670 ;
      RECT 53.4950 80.8100 54.9960 82.3540 ;
      RECT 54.0960 77.8180 54.9960 78.3640 ;
      RECT 0.0000 0.0000 19.9860 0.9000 ;
      RECT 0.0000 61.7520 54.9960 67.3980 ;
      RECT 0.9000 61.7000 54.9960 67.3980 ;
      RECT 0.9000 58.6270 54.0960 67.3980 ;
      RECT 0.9000 61.7000 54.9960 61.7520 ;
      RECT 0.9000 58.6270 54.0960 61.7000 ;
      RECT 0.0000 67.3980 54.0960 67.4490 ;
      RECT 0.0000 61.7520 54.0960 67.4490 ;
      RECT 0.9000 67.4490 54.0960 70.5190 ;
      RECT 0.9000 61.7520 54.0960 70.5190 ;
      RECT 0.0000 83.9540 54.9960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 90.2530 ;
      RECT 0.0000 83.9030 54.0960 83.9540 ;
      RECT 0.9000 82.3540 54.0960 83.9030 ;
      RECT 0.0000 58.5810 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.0960 58.6270 ;
      RECT 0.0000 26.8660 54.9960 58.5810 ;
      RECT 0.9000 26.8660 54.0960 61.7000 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 58.5810 ;
      RECT 0.9000 26.8610 54.9960 26.8660 ;
      RECT 0.9000 25.2660 54.0960 26.8610 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.9000 28.1480 9.1540 ;
      RECT 0.0000 0.0000 19.9860 9.1540 ;
      RECT 0.0000 0.9000 28.1480 0.9010 ;
      RECT 0.9000 9.1560 54.0960 10.7540 ;
      RECT 0.0000 25.2610 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.0960 25.2660 ;
      RECT 0.0000 18.3290 54.9960 25.2610 ;
      RECT 0.0000 16.1630 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.0960 16.1680 ;
      RECT 0.0000 10.7560 54.9960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 16.1630 ;
      RECT 0.0000 10.7540 54.0960 10.7560 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.3290 54.0960 26.8610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 25.2610 ;
      RECT 0.9000 10.7560 54.0960 25.2610 ;
      RECT 0.9000 10.7560 54.0960 25.2610 ;
      RECT 0.9000 10.7560 54.0960 25.2610 ;
      RECT 0.9000 18.2330 54.9960 18.3290 ;
      RECT 0.9000 16.1680 54.0960 18.2330 ;
      RECT 0.0000 0.9010 54.9960 9.1540 ;
      RECT 0.9000 9.1540 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 0.9000 0.9010 54.9960 9.1560 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 9.1540 ;
      RECT 29.7480 0.9000 54.9960 0.9010 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 9.1540 ;
      RECT 35.0180 0.0000 54.9960 0.9000 ;
      RECT 0.9000 79.1510 54.0960 90.2530 ;
      RECT 0.9000 79.1510 54.0960 90.2530 ;
      RECT 0.9000 80.8100 54.0960 83.9540 ;
      RECT 0.9000 79.1510 54.0960 83.9540 ;
      RECT 0.9000 79.1510 54.0960 83.9540 ;
      RECT 0.9000 80.8100 54.0960 83.9030 ;
      RECT 0.9000 80.8100 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 80.7510 54.0960 83.9030 ;
      RECT 0.9000 82.3030 54.0960 82.3540 ;
      RECT 0.9000 79.1510 54.0960 82.3540 ;
      RECT 0.9000 79.1510 54.0960 82.3540 ;
      RECT 0.9000 80.8100 54.0960 82.3030 ;
      RECT 0.0000 70.5710 54.9960 76.2180 ;
      RECT 0.9000 70.5190 54.9960 70.5710 ;
      RECT 0.9000 67.4490 54.0960 70.5710 ;
      RECT 0.9000 76.2670 54.0960 90.2530 ;
      RECT 0.9000 76.2670 54.0960 90.2530 ;
      RECT 0.9000 76.2670 54.0960 83.9540 ;
      RECT 0.9000 76.2670 54.0960 82.3540 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 82.3030 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.8100 ;
      RECT 0.9000 76.2670 54.0960 80.7510 ;
      RECT 0.9000 78.3640 54.0960 79.1510 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 54.9960 90.2530 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 54.9960 90.2530 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 54.9960 90.2530 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 54.9960 90.2530 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 54.9960 90.2530 ;
  END
END SRAMLP2RW64x4

MACRO SRAMLP2RW64x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 67.056 BY 92.317 ;
  SYMMETRY X Y R90 ;

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.8700 0.0010 42.0700 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.8700 0.0010 42.0700 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.8700 0.0010 42.0700 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.8700 0.0010 42.0700 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.8700 0.0010 42.0700 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.6060 0.0000 44.8060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.6060 0.0010 44.8060 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.6060 0.0010 44.8060 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.6060 0.0010 44.8060 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.6060 0.0010 44.8060 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.2380 0.0010 43.4380 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.2380 0.0010 43.4380 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.2380 0.0010 43.4380 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.2380 0.0010 43.4380 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.2380 0.0010 43.4380 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.2770 0.0000 45.4770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.2770 0.0010 45.4770 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.2770 0.0010 45.4770 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.2770 0.0010 45.4770 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.2770 0.0010 45.4770 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.2600 0.0010 33.4600 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.2600 0.0010 33.4600 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.2600 0.0010 33.4600 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.2600 0.0010 33.4600 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.2600 0.0010 33.4600 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.9310 0.0010 34.1310 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.9310 0.0010 34.1310 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.9310 0.0010 34.1310 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.9310 0.0010 34.1310 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.9310 0.0010 34.1310 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 81.1700 67.0560 81.3700 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 81.1700 67.0560 81.3700 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 81.1700 67.0560 81.3700 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 81.1700 67.0560 81.3700 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 81.1700 67.0560 81.3700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAGATEAREA 0.0792 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 4.116344 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.116344 LAYER M3 ;
    ANTENNAMAXAREACAR 54.93026 LAYER M3 ;
    ANTENNAGATEAREA 0.0792 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 56.81548 LAYER M4 ;
    ANTENNAGATEAREA 0.0792 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 58.70057 LAYER M5 ;
    ANTENNAGATEAREA 0.0792 LAYER M6 ;
    ANTENNAGATEAREA 0.0792 LAYER M7 ;
    ANTENNAGATEAREA 0.0792 LAYER M8 ;
    ANTENNAGATEAREA 0.0792 LAYER M9 ;
    ANTENNAGATEAREA 0.0792 LAYER MRDL ;
  END SD

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 85.1970 67.0560 85.3970 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 85.1970 67.0560 85.3970 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 85.1970 67.0560 85.3970 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 85.1970 67.0560 85.3970 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 85.1970 67.0560 85.3970 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.202265 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.202265 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.938872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.938872 LAYER M2 ;
    ANTENNAMAXAREACAR 20.81647 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.42173 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 30.46409 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.50626 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 82.0530 67.0560 82.2530 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 82.0530 67.0560 82.2530 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 82.0530 67.0560 82.2530 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 82.0530 67.0560 82.2530 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 82.0530 67.0560 82.2530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.208108 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.208108 LAYER M2 ;
    ANTENNAMAXAREACAR 11.2157 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 3.686098 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.686098 LAYER M3 ;
    ANTENNAMAXAREACAR 82.44756 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 95.32571 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 98.60004 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS1

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 82.0320 0.2000 82.2320 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 82.0320 0.2000 82.2320 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 82.0320 0.2000 82.2320 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 82.0320 0.2000 82.2320 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 82.0320 0.2000 82.2320 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16318 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16318 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.239388 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.239388 LAYER M2 ;
    ANTENNAMAXAREACAR 12.68426 LAYER M2 ;
    ANTENNAGATEAREA 0.0456 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.233183 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.233183 LAYER M3 ;
    ANTENNAMAXAREACAR 28.36307 LAYER M3 ;
    ANTENNAGATEAREA 0.0456 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 43.04958 LAYER M4 ;
    ANTENNAGATEAREA 0.0456 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 46.37131 LAYER M5 ;
    ANTENNAGATEAREA 0.0456 LAYER M6 ;
    ANTENNAGATEAREA 0.0456 LAYER M7 ;
    ANTENNAGATEAREA 0.0456 LAYER M8 ;
    ANTENNAGATEAREA 0.0456 LAYER M9 ;
    ANTENNAGATEAREA 0.0456 LAYER MRDL ;
  END DS2

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 85.1840 0.2000 85.3840 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 85.1840 0.2000 85.3840 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 85.1840 0.2000 85.3840 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 85.1840 0.2000 85.3840 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 85.1840 0.2000 85.3840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.230665 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.230665 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.938872 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.938872 LAYER M2 ;
    ANTENNAMAXAREACAR 20.81647 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 28.19762 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.23994 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.28206 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.3910 0.0000 21.5910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.3910 0.0000 21.5910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.3910 0.0000 21.5910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.3910 0.0000 21.5910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.3910 0.0000 21.5910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.90238 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.90238 LAYER M2 ;
    ANTENNAMAXAREACAR 7.258762 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.315466 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.372101 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.42867 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.7670 0.0000 45.9670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.7670 0.0000 45.9670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.7670 0.0000 45.9670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.7670 0.0000 45.9670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.7670 0.0000 45.9670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.9076 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9076 LAYER M2 ;
    ANTENNAMAXAREACAR 7.295164 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.351866 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.408497 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.46506 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB1

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 9.8570 67.0560 10.0570 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 9.8570 67.0560 10.0570 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 9.8570 67.0560 10.0570 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 9.8570 67.0560 10.0570 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 9.8570 67.0560 10.0570 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.59754 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.59754 LAYER M2 ;
    ANTENNAMAXAREACAR 11.9729 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 13.00976 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.04654 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.08326 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8560 0.2000 10.0560 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8560 0.2000 10.0560 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8560 0.2000 10.0560 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8560 0.2000 10.0560 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8560 0.2000 10.0560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.61614 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.61614 LAYER M2 ;
    ANTENNAMAXAREACAR 12.10021 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 13.13706 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.17384 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 15.21055 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.0300 0.0010 35.2300 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.0300 0.0010 35.2300 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.0300 0.0010 35.2300 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.0300 0.0010 35.2300 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.0300 0.0010 35.2300 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.3980 0.0010 36.5980 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.3980 0.0010 36.5980 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.3980 0.0010 36.5980 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.3980 0.0010 36.5980 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.3980 0.0010 36.5980 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.7230 0.0010 25.9230 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.7230 0.0010 25.9230 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.7230 0.0010 25.9230 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.7230 0.0010 25.9230 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.7230 0.0010 25.9230 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.4200 0.0010 26.6200 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.4200 0.0010 26.6200 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.4200 0.0010 26.6200 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.4200 0.0010 26.6200 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.4200 0.0010 26.6200 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.7880 0.0010 27.9880 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.7880 0.0010 27.9880 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.7880 0.0010 27.9880 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.7880 0.0010 27.9880 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.7880 0.0010 27.9880 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.8270 0.0010 30.0270 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.8270 0.0010 30.0270 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.8270 0.0010 30.0270 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.8270 0.0010 30.0270 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.8270 0.0010 30.0270 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.4590 0.0010 28.6590 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.4590 0.0010 28.6590 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.4590 0.0010 28.6590 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.4590 0.0010 28.6590 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.4590 0.0010 28.6590 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.1560 0.0010 29.3560 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.1560 0.0010 29.3560 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.1560 0.0010 29.3560 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.1560 0.0010 29.3560 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.1560 0.0010 29.3560 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.5240 0.0010 30.7240 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.5240 0.0010 30.7240 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.5240 0.0010 30.7240 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.5240 0.0010 30.7240 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.5240 0.0010 30.7240 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.7660 0.0010 37.9660 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.7660 0.0010 37.9660 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.7660 0.0010 37.9660 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.7660 0.0010 37.9660 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.7660 0.0010 37.9660 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.5630 0.0010 32.7630 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.5630 0.0010 32.7630 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.5630 0.0010 32.7630 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.5630 0.0010 32.7630 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.5630 0.0010 32.7630 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.8920 0.0010 32.0920 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.8920 0.0010 32.0920 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.8920 0.0010 32.0920 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.8920 0.0010 32.0920 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.8920 0.0010 32.0920 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.7010 0.0010 35.9010 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.7010 0.0010 35.9010 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.7010 0.0010 35.9010 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.7010 0.0010 35.9010 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.7010 0.0010 35.9010 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.4370 0.0010 38.6370 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.4370 0.0010 38.6370 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.4370 0.0010 38.6370 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.4370 0.0010 38.6370 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.4370 0.0010 38.6370 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.1950 0.0010 31.3950 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.1950 0.0010 31.3950 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.1950 0.0010 31.3950 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.1950 0.0010 31.3950 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.1950 0.0010 31.3950 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.1340 0.0010 39.3340 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.1340 0.0010 39.3340 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.1340 0.0010 39.3340 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.1340 0.0010 39.3340 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.1340 0.0010 39.3340 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.1730 0.0010 41.3730 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.1730 0.0010 41.3730 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.1730 0.0010 41.3730 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.1730 0.0010 41.3730 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.1730 0.0010 41.3730 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.8050 0.0010 40.0050 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.8050 0.0010 40.0050 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.8050 0.0010 40.0050 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.8050 0.0010 40.0050 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.8050 0.0010 40.0050 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.5410 0.0010 42.7410 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.5410 0.0010 42.7410 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.5410 0.0010 42.7410 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.5410 0.0010 42.7410 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.5410 0.0010 42.7410 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5020 0.0010 40.7020 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5020 0.0010 40.7020 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5020 0.0010 40.7020 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5020 0.0010 40.7020 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5020 0.0010 40.7020 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.9090 0.0010 44.1090 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.9090 0.0010 44.1090 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.9090 0.0010 44.1090 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.9090 0.0010 44.1090 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.9090 0.0010 44.1090 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.1250 0.2000 28.3250 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 28.1250 0.2000 28.3250 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 28.1250 0.2000 28.3250 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 28.1250 0.2000 28.3250 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 28.1250 0.2000 28.3250 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.182128 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.182128 LAYER M4 ;
    ANTENNAMAXAREACAR 59.94311 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 67.15821 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[5]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.0690 0.0010 37.2690 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.0690 0.0010 37.2690 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.0690 0.0010 37.2690 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.0690 0.0010 37.2690 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.0690 0.0010 37.2690 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8690 0.2000 17.0690 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8690 0.2000 17.0690 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8690 0.2000 17.0690 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8690 0.2000 17.0690 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8690 0.2000 17.0690 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.474112 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.474112 LAYER M4 ;
    ANTENNAMAXAREACAR 15.26801 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 19.40908 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4300 0.2000 17.6300 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4300 0.2000 17.6300 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4300 0.2000 17.6300 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4300 0.2000 17.6300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4300 0.2000 17.6300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.358 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.358 LAYER M4 ;
    ANTENNAMAXAREACAR 13.89914 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.33097 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 79.0780 67.0560 79.2780 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 79.0780 67.0560 79.2780 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 79.0780 67.0560 79.2780 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 79.0780 67.0560 79.2780 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 79.0780 67.0560 79.2780 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.940008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.940008 LAYER M3 ;
    ANTENNAMAXAREACAR 27.47615 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 31.56175 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 35.64707 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[0]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 70.2580 67.0560 70.4580 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 70.2580 67.0560 70.4580 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 70.2580 67.0560 70.4580 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 70.2580 67.0560 70.4580 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 70.2580 67.0560 70.4580 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.941408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941408 LAYER M3 ;
    ANTENNAMAXAREACAR 27.5144 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.65467 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.79465 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 71.7790 67.0560 71.9790 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 71.7790 67.0560 71.9790 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 71.7790 67.0560 71.9790 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 71.7790 67.0560 71.9790 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 71.7790 67.0560 71.9790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.940008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.940008 LAYER M3 ;
    ANTENNAMAXAREACAR 27.47615 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M4 ;
    ANTENNAMAXAREACAR 31.56175 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1496 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1496 LAYER M5 ;
    ANTENNAMAXAREACAR 35.64707 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[1]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 61.4390 67.0560 61.6390 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 61.4390 67.0560 61.6390 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 61.4390 67.0560 61.6390 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 61.4390 67.0560 61.6390 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 61.4390 67.0560 61.6390 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.941408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941408 LAYER M3 ;
    ANTENNAMAXAREACAR 27.5144 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.65467 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.79465 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[4]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 62.9600 67.0560 63.1600 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 62.9600 67.0560 63.1600 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 62.9600 67.0560 63.1600 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 62.9600 67.0560 63.1600 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 62.9600 67.0560 63.1600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.941408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941408 LAYER M3 ;
    ANTENNAMAXAREACAR 27.5144 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.65467 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.79465 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[3]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 28.1210 67.0560 28.3210 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 28.1210 67.0560 28.3210 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 28.1210 67.0560 28.3210 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 28.1210 67.0560 28.3210 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 28.1210 67.0560 28.3210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.163491 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.163491 LAYER M4 ;
    ANTENNAMAXAREACAR 58.89658 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 66.11175 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[5]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 16.8650 67.0560 17.0650 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 16.8650 67.0560 17.0650 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 16.8650 67.0560 17.0650 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 16.8650 67.0560 17.0650 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 16.8650 67.0560 17.0650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.452569 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.452569 LAYER M4 ;
    ANTENNAMAXAREACAR 14.29994 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.44107 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8560 17.3340 67.0560 17.5340 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8560 17.3340 67.0560 17.5340 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8560 17.3340 67.0560 17.5340 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8560 17.3340 67.0560 17.5340 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8560 17.3340 67.0560 17.5340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.32974 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.32974 LAYER M4 ;
    ANTENNAMAXAREACAR 13.42818 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.86005 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 16.2220 92.0160 16.5220 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1220 92.0160 17.4220 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6210 92.0160 3.9220 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.5210 92.0160 4.8210 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.1210 92.0160 62.4200 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.0210 92.0160 63.3200 92.3160 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 164.4285 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 164.4285 LAYER M5 ;
  END VDDL

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 79.1270 0.2000 79.3270 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 79.1270 0.2000 79.3270 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 79.1270 0.2000 79.3270 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 79.1270 0.2000 79.3270 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 79.1270 0.2000 79.3270 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.960008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.960008 LAYER M3 ;
    ANTENNAMAXAREACAR 28.0226 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 32.16283 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.30279 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.3550 0.0010 24.5550 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.3550 0.0010 24.5550 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.3550 0.0010 24.5550 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.3550 0.0010 24.5550 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.3550 0.0010 24.5550 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.6840 0.0010 23.8840 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.6840 0.0010 23.8840 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.6840 0.0010 23.8840 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.6840 0.0010 23.8840 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.6840 0.0010 23.8840 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.0520 0.0010 25.2520 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.0520 0.0010 25.2520 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.0520 0.0010 25.2520 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.0520 0.0010 25.2520 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.0520 0.0010 25.2520 0.2010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.285988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285988 LAYER M3 ;
    ANTENNAMAXAREACAR 62.48578 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.70071 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.91516 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.0910 0.0010 27.2910 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.0910 0.0010 27.2910 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.0910 0.0010 27.2910 0.2010 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.0910 0.0010 27.2910 0.2010 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.0910 0.0010 27.2910 0.2010 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26188 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 71.8280 0.2000 72.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 71.8280 0.2000 72.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 71.8280 0.2000 72.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 71.8280 0.2000 72.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 71.8280 0.2000 72.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.960008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.960008 LAYER M3 ;
    ANTENNAMAXAREACAR 28.0226 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 32.16283 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.30279 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 70.3100 0.2000 70.5100 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 70.3100 0.2000 70.5100 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 70.3100 0.2000 70.5100 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 70.3100 0.2000 70.5100 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 70.3100 0.2000 70.5100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.960008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.960008 LAYER M3 ;
    ANTENNAMAXAREACAR 28.0226 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 32.16283 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.30279 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 61.4870 0.2000 61.6870 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 61.4870 0.2000 61.6870 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 61.4870 0.2000 61.6870 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 61.4870 0.2000 61.6870 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 61.4870 0.2000 61.6870 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.960008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.960008 LAYER M3 ;
    ANTENNAMAXAREACAR 28.0226 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 32.16283 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.30279 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[4]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 63.0120 0.2000 63.2120 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 63.0120 0.2000 63.2120 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 63.0120 0.2000 63.2120 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 63.0120 0.2000 63.2120 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 63.0120 0.2000 63.2120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.960728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.960728 LAYER M3 ;
    ANTENNAMAXAREACAR 28.06524 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 32.20546 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 36.34541 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[3]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 1.8200 92.0160 2.1190 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7220 92.0160 3.0210 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6210 92.0160 12.9220 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7210 92.0160 12.0220 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.3220 92.0160 51.6220 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.8200 92.0160 65.1190 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.4210 92.0160 50.7210 92.3160 ;
    END
    ANTENNADIFFAREA 10.95167 LAYER M5 ;
    ANTENNADIFFAREA 10.95167 LAYER M6 ;
    ANTENNADIFFAREA 10.95167 LAYER M7 ;
    ANTENNADIFFAREA 10.95167 LAYER M8 ;
    ANTENNADIFFAREA 10.95167 LAYER M9 ;
    ANTENNADIFFAREA 10.95167 LAYER MRDL ;
    ANTENNAGATEAREA 1.5408 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 629.511 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 629.511 LAYER M5 ;
    ANTENNAMAXAREACAR 447.3804 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 164.4288 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 164.4288 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 22.0710 92.0160 22.3710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.4700 92.0160 63.7700 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.2700 92.0160 65.5700 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.7710 92.0160 52.0710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.5720 92.0160 53.8720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.1720 92.0160 57.4720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.7720 92.0160 61.0720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.5710 92.0160 62.8710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.6710 92.0160 61.9710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.8710 92.0160 60.1710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.9710 92.0160 59.2710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.0710 92.0160 58.3710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.2710 92.0160 56.5710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.3710 92.0160 55.6710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.4710 92.0160 54.7710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.6710 92.0160 52.9710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.6710 92.0160 43.9710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.7710 92.0160 43.0710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.0720 92.0160 49.3720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.3720 92.0160 46.6730 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.4710 92.0160 45.7700 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.8720 92.0160 42.1730 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.5720 92.0160 44.8720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.9710 92.0160 50.2700 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.1710 92.0160 48.4710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.2710 92.0160 47.5710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.5720 92.0160 35.8710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.7720 92.0160 34.0720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.9710 92.0160 41.2700 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.0720 92.0160 40.3720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.1710 92.0160 39.4710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.2710 92.0160 38.5710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.6720 92.0160 34.9710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.1720 92.0160 30.4710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.4710 92.0160 36.7720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.0720 92.0160 31.3710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.4720 92.0160 27.7720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.2720 92.0160 29.5720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.6710 92.0160 16.9710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.9710 92.0160 23.2720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.4710 92.0160 9.7720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.8710 92.0160 15.1710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.6710 92.0160 25.9720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.8720 92.0160 24.1720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1720 92.0160 12.4710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.1720 92.0160 3.4720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2710 92.0160 2.5710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.9720 92.0160 14.2720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.5720 92.0160 8.8710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.7720 92.0160 16.0710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.3710 92.0160 10.6720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.0710 92.0160 4.3710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.2720 92.0160 11.5720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.0710 92.0160 13.3710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.3710 92.0160 19.6720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.7720 92.0160 7.0720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.1720 92.0160 21.4720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8710 92.0160 6.1720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.2720 92.0160 20.5720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.3710 92.0160 28.6710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.5710 92.0160 17.8720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.6720 92.0160 7.9710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4710 92.0160 18.7720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.8710 92.0160 33.1720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.9710 92.0160 32.2720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9710 92.0160 5.2720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.5710 92.0160 26.8710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.7720 92.0160 25.0710 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.3710 92.0160 37.6720 92.3160 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.3710 92.0160 64.6710 92.3160 ;
    END
    ANTENNADIFFAREA 151.4734 LAYER M5 ;
    ANTENNADIFFAREA 151.4734 LAYER M6 ;
    ANTENNADIFFAREA 151.4734 LAYER M7 ;
    ANTENNADIFFAREA 151.4734 LAYER M8 ;
    ANTENNADIFFAREA 151.4734 LAYER M9 ;
    ANTENNADIFFAREA 151.4734 LAYER MRDL ;
    ANTENNAGATEAREA 5.49 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1939.135 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 1939.135 LAYER M5 ;
    ANTENNAMAXAREACAR 439.5299 LAYER M5 ;
    ANTENNAGATEAREA 5.49 LAYER M6 ;
    ANTENNAGATEAREA 5.49 LAYER M7 ;
    ANTENNAGATEAREA 5.49 LAYER M8 ;
    ANTENNAGATEAREA 5.49 LAYER M9 ;
    ANTENNAGATEAREA 5.49 LAYER MRDL ;
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.8000 28.9210 67.0560 60.8390 ;
      RECT 0.8000 28.9210 67.0560 60.8390 ;
      RECT 0.8000 28.9210 67.0560 60.8390 ;
      RECT 0.8000 28.9210 67.0560 28.9250 ;
      RECT 0.8000 82.8530 66.2560 85.9970 ;
      RECT 0.0000 72.6280 67.0560 78.4780 ;
      RECT 0.0000 63.8120 67.0560 69.6580 ;
      RECT 0.8000 69.7100 66.2560 72.5790 ;
      RECT 0.8000 60.8870 66.2560 69.6580 ;
      RECT 0.8000 60.8870 66.2560 69.6580 ;
      RECT 0.8000 60.8870 66.2560 69.6580 ;
      RECT 0.8000 60.8870 66.2560 69.6580 ;
      RECT 0.8000 60.8870 66.2560 69.6580 ;
      RECT 0.8000 60.8870 66.2560 69.6580 ;
      RECT 0.8000 60.8390 66.2560 69.6580 ;
      RECT 0.8000 60.8390 66.2560 69.6580 ;
      RECT 0.8000 60.8390 66.2560 69.6580 ;
      RECT 0.8000 78.5270 66.2560 85.9840 ;
      RECT 0.8000 78.5270 66.2560 82.8320 ;
      RECT 0.8000 78.5270 66.2560 82.8320 ;
      RECT 0.8000 78.5270 66.2560 82.8320 ;
      RECT 22.1910 0.0000 23.0840 0.8000 ;
      RECT 0.0000 79.9270 1.5010 81.4320 ;
      RECT 0.0000 66.7090 66.2560 69.7100 ;
      RECT 0.0000 82.8320 1.5010 84.5840 ;
      RECT 0.0000 60.8390 3.0010 60.8870 ;
      RECT 66.2560 79.8780 67.0560 80.5700 ;
      RECT 64.0550 63.7600 67.0560 63.8120 ;
      RECT 65.5550 82.8530 67.0560 84.5970 ;
      RECT 66.2560 71.1590 67.0560 71.1790 ;
      RECT 0.8000 71.0580 67.0560 71.1100 ;
      RECT 0.8000 69.7100 66.2560 71.0580 ;
      RECT 0.0000 75.5800 66.2560 78.5270 ;
      RECT 0.0000 75.5260 67.0560 75.5800 ;
      RECT 0.8000 72.5790 67.0560 75.5260 ;
      RECT 0.0000 71.1100 67.0560 71.1590 ;
      RECT 0.0000 62.2870 0.8000 62.4120 ;
      RECT 66.2560 62.2390 67.0560 62.3600 ;
      RECT 0.0000 71.1590 0.8000 71.2280 ;
      RECT 0.0000 0.0000 20.7910 0.8000 ;
      RECT 0.0000 10.6570 67.0560 16.2650 ;
      RECT 0.0000 0.8000 23.0840 0.8010 ;
      RECT 0.0000 0.0000 20.7910 9.2560 ;
      RECT 0.0000 0.0000 20.7910 9.2560 ;
      RECT 0.0000 0.8000 23.0840 9.2560 ;
      RECT 0.0000 0.8000 23.0840 9.2560 ;
      RECT 0.0000 85.9970 67.0560 92.3170 ;
      RECT 0.0000 85.9840 66.2560 85.9970 ;
      RECT 0.0000 16.2650 66.2560 16.2690 ;
      RECT 0.0000 10.6570 66.2560 16.2690 ;
      RECT 0.0000 10.6570 66.2560 16.2690 ;
      RECT 0.0000 10.6570 66.2560 16.2690 ;
      RECT 0.8000 16.2690 66.2560 18.1340 ;
      RECT 0.0000 10.6560 66.2560 16.2650 ;
      RECT 0.0000 10.6560 66.2560 16.2650 ;
      RECT 0.0000 10.6560 66.2560 16.2650 ;
      RECT 0.0000 10.6560 66.2560 10.6570 ;
      RECT 0.8000 9.2570 66.2560 10.6560 ;
      RECT 0.0000 27.5210 66.2560 27.5250 ;
      RECT 0.0000 18.2300 66.2560 27.5250 ;
      RECT 0.0000 18.2300 66.2560 27.5250 ;
      RECT 0.0000 18.2300 66.2560 27.5250 ;
      RECT 0.0000 18.2300 67.0560 27.5210 ;
      RECT 0.8000 18.1340 67.0560 27.5210 ;
      RECT 0.8000 18.1340 67.0560 27.5210 ;
      RECT 0.8000 18.1340 67.0560 27.5210 ;
      RECT 0.8000 10.6570 66.2560 27.5210 ;
      RECT 0.8000 10.6570 66.2560 27.5210 ;
      RECT 0.8000 10.6570 66.2560 27.5210 ;
      RECT 0.8000 18.1340 67.0560 18.2300 ;
      RECT 0.8000 27.5250 66.2560 28.9210 ;
      RECT 0.8000 18.2300 66.2560 28.9210 ;
      RECT 0.8000 18.2300 66.2560 28.9210 ;
      RECT 0.8000 18.2300 66.2560 28.9210 ;
      RECT 0.0000 0.8010 67.0560 9.2560 ;
      RECT 0.8000 9.2560 67.0560 9.2570 ;
      RECT 0.8000 0.8010 67.0560 9.2570 ;
      RECT 0.8000 0.8010 67.0560 9.2570 ;
      RECT 0.8000 0.8010 67.0560 9.2570 ;
      RECT 46.0770 0.8000 67.0560 9.2560 ;
      RECT 46.0770 0.8000 67.0560 9.2560 ;
      RECT 46.0770 0.8000 67.0560 0.8010 ;
      RECT 46.5670 0.0000 67.0560 9.2560 ;
      RECT 46.5670 0.0000 67.0560 9.2560 ;
      RECT 46.5670 0.0000 67.0560 0.8000 ;
      RECT 0.0000 28.9250 67.0560 60.8390 ;
      RECT 0.8000 60.8870 66.2560 63.7600 ;
    LAYER PO ;
      RECT 0.0000 0.0000 67.0560 92.3170 ;
    LAYER M2 ;
      RECT 0.0000 16.1650 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 67.0560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 10.7570 ;
      RECT 0.9000 16.1690 66.1560 18.2340 ;
      RECT 0.0000 27.4210 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 18.3300 ;
      RECT 0.0000 69.5580 66.1560 69.6100 ;
      RECT 0.0000 63.9120 66.1560 69.6100 ;
      RECT 0.0000 63.9120 67.0560 69.5580 ;
      RECT 0.9000 63.9120 66.1560 72.6790 ;
      RECT 0.9000 63.8600 67.0560 69.5580 ;
      RECT 0.9000 60.7870 66.1560 69.5580 ;
      RECT 0.9000 63.8600 67.0560 63.9120 ;
      RECT 0.9000 60.7870 66.1560 63.8600 ;
      RECT 0.0000 60.7390 66.1560 60.7870 ;
      RECT 0.0000 29.0250 66.1560 60.7870 ;
      RECT 0.0000 29.0250 67.0560 60.7390 ;
      RECT 0.9000 29.0250 66.1560 63.8600 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 29.0250 ;
      RECT 0.9000 27.4250 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.0000 0.9010 67.0560 9.1560 ;
      RECT 0.9000 9.1560 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 46.1770 0.9000 67.0560 9.1560 ;
      RECT 46.1770 0.9000 67.0560 9.1560 ;
      RECT 46.1770 0.9000 67.0560 0.9010 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 0.9000 ;
      RECT 0.0000 72.7280 67.0560 78.3780 ;
      RECT 0.9000 72.6790 67.0560 72.7280 ;
      RECT 0.9000 69.6100 66.1560 72.7280 ;
      RECT 0.9000 82.9530 66.1560 86.0970 ;
      RECT 0.9000 78.4270 66.1560 86.0840 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 22.2910 0.0000 22.9840 0.9000 ;
      RECT 0.0000 75.4260 66.1560 78.4270 ;
      RECT 0.0000 82.9320 1.5010 84.4840 ;
      RECT 66.1560 79.9780 67.0560 80.4700 ;
      RECT 65.5550 82.9530 67.0560 84.4970 ;
      RECT 0.0000 80.0270 0.9000 81.3320 ;
      RECT 0.0000 0.0000 20.6910 0.9000 ;
      RECT 0.0000 0.9000 22.9840 0.9010 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.9000 9.1570 66.1560 10.7560 ;
      RECT 0.9000 69.6100 66.1560 72.6790 ;
      RECT 0.0000 86.0970 67.0560 92.3170 ;
      RECT 0.0000 86.0840 66.1560 86.0970 ;
    LAYER M4 ;
      RECT 0.9000 60.7870 66.1560 69.5580 ;
      RECT 0.9000 63.8600 67.0560 63.9120 ;
      RECT 0.9000 60.7870 66.1560 63.8600 ;
      RECT 0.0000 60.7390 66.1560 60.7870 ;
      RECT 0.0000 29.0250 66.1560 60.7870 ;
      RECT 0.0000 29.0250 67.0560 60.7390 ;
      RECT 0.9000 29.0250 66.1560 63.8600 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 29.0250 ;
      RECT 0.9000 27.4250 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.0000 0.9010 67.0560 9.1560 ;
      RECT 0.9000 9.1560 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 46.1770 0.9000 67.0560 9.1560 ;
      RECT 46.1770 0.9000 67.0560 9.1560 ;
      RECT 46.1770 0.9000 67.0560 0.9010 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 0.9000 ;
      RECT 0.0000 72.7280 67.0560 78.3780 ;
      RECT 0.9000 72.6790 67.0560 72.7280 ;
      RECT 0.9000 69.6100 66.1560 72.7280 ;
      RECT 0.9000 82.9530 66.1560 86.0970 ;
      RECT 0.9000 78.4270 66.1560 86.0840 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 22.2910 0.0000 22.9840 0.9000 ;
      RECT 0.0000 80.0270 0.9000 81.3320 ;
      RECT 0.0000 82.9320 1.5010 84.4840 ;
      RECT 0.0000 75.4260 66.1560 78.4270 ;
      RECT 65.5550 82.9530 67.0560 84.4970 ;
      RECT 66.1560 79.9780 67.0560 80.4700 ;
      RECT 0.0000 0.0000 20.6910 0.9000 ;
      RECT 0.0000 0.9000 22.9840 0.9010 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.9000 9.1570 66.1560 10.7560 ;
      RECT 0.9000 69.6100 66.1560 72.6790 ;
      RECT 0.0000 86.0970 67.0560 92.3170 ;
      RECT 0.0000 86.0840 66.1560 86.0970 ;
      RECT 0.0000 16.1650 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 67.0560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 10.7570 ;
      RECT 0.9000 16.1690 66.1560 18.2340 ;
      RECT 0.0000 27.4210 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 18.3300 ;
      RECT 0.0000 69.5580 66.1560 69.6100 ;
      RECT 0.0000 63.9120 66.1560 69.6100 ;
      RECT 0.0000 63.9120 67.0560 69.5580 ;
      RECT 0.9000 63.9120 66.1560 72.6790 ;
      RECT 0.9000 63.8600 67.0560 69.5580 ;
    LAYER M3 ;
      RECT 22.2910 0.0000 22.9840 0.9000 ;
      RECT 0.0000 80.0270 0.9000 81.3320 ;
      RECT 0.0000 82.9320 1.5010 84.4840 ;
      RECT 0.0000 75.4260 66.1560 78.4270 ;
      RECT 65.5550 82.9530 67.0560 84.4970 ;
      RECT 66.1560 79.9780 67.0560 80.4700 ;
      RECT 0.0000 0.0000 20.6910 0.9000 ;
      RECT 0.0000 0.9000 22.9840 0.9010 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.9000 9.1570 66.1560 10.7560 ;
      RECT 0.9000 69.6100 66.1560 72.6790 ;
      RECT 0.0000 86.0970 67.0560 92.3170 ;
      RECT 0.0000 86.0840 66.1560 86.0970 ;
      RECT 0.0000 16.1650 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 67.0560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 10.7570 ;
      RECT 0.9000 16.1690 66.1560 18.2340 ;
      RECT 0.0000 27.4210 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 18.3300 ;
      RECT 0.0000 69.5580 66.1560 69.6100 ;
      RECT 0.0000 63.9120 66.1560 69.6100 ;
      RECT 0.0000 63.9120 67.0560 69.5580 ;
      RECT 0.9000 63.9120 66.1560 72.6790 ;
      RECT 0.9000 63.8600 67.0560 69.5580 ;
      RECT 0.9000 60.7870 66.1560 69.5580 ;
      RECT 0.9000 63.8600 67.0560 63.9120 ;
      RECT 0.9000 60.7870 66.1560 63.8600 ;
      RECT 0.0000 60.7390 66.1560 60.7870 ;
      RECT 0.0000 29.0250 66.1560 60.7870 ;
      RECT 0.0000 29.0250 67.0560 60.7390 ;
      RECT 0.9000 29.0250 66.1560 63.8600 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 29.0250 ;
      RECT 0.9000 27.4250 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.0000 0.9010 67.0560 9.1560 ;
      RECT 0.9000 9.1560 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 46.1770 0.9000 67.0560 9.1560 ;
      RECT 46.1770 0.9000 67.0560 9.1560 ;
      RECT 46.1770 0.9000 67.0560 0.9010 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 0.9000 ;
      RECT 0.0000 72.7280 67.0560 78.3780 ;
      RECT 0.9000 72.6790 67.0560 72.7280 ;
      RECT 0.9000 69.6100 66.1560 72.7280 ;
      RECT 0.9000 82.9530 66.1560 86.0970 ;
      RECT 0.9000 78.4270 66.1560 86.0840 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 67.0560 92.3170 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 67.0560 92.3170 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 67.0560 92.3170 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 67.0560 92.3170 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 67.0560 92.3170 ;
    LAYER M5 ;
      RECT 0.0000 91.3160 1.1200 92.3170 ;
      RECT 22.2910 0.0000 22.9840 0.9000 ;
      RECT 66.2700 91.3160 67.0560 92.3170 ;
      RECT 0.0000 80.0270 0.9000 81.3320 ;
      RECT 0.0000 75.4260 66.1560 78.4270 ;
      RECT 0.0000 82.9320 1.5010 84.4840 ;
      RECT 65.5550 82.9530 67.0560 84.4970 ;
      RECT 66.1560 79.9780 67.0560 80.4700 ;
      RECT 0.0000 0.0000 20.6910 0.9000 ;
      RECT 0.0000 0.9000 22.9840 0.9010 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.0000 20.6910 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.0000 0.9000 22.9840 9.1560 ;
      RECT 0.9000 9.1570 66.1560 10.7560 ;
      RECT 0.9000 69.6100 66.1560 72.6790 ;
      RECT 0.0000 86.0970 67.0560 91.3160 ;
      RECT 0.0000 86.0840 66.1560 86.0970 ;
      RECT 0.0000 16.1650 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 66.1560 16.1690 ;
      RECT 0.0000 10.7570 67.0560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 16.1650 ;
      RECT 0.0000 10.7560 66.1560 10.7570 ;
      RECT 0.9000 16.1690 66.1560 18.2340 ;
      RECT 0.0000 27.4210 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 66.1560 27.4250 ;
      RECT 0.0000 18.3300 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 10.7570 66.1560 27.4210 ;
      RECT 0.9000 18.2340 67.0560 18.3300 ;
      RECT 0.0000 69.5580 66.1560 69.6100 ;
      RECT 0.0000 63.9120 66.1560 69.6100 ;
      RECT 0.0000 63.9120 67.0560 69.5580 ;
      RECT 0.9000 63.9120 66.1560 72.6790 ;
      RECT 0.9000 63.8600 67.0560 69.5580 ;
      RECT 0.9000 60.7870 66.1560 69.5580 ;
      RECT 0.9000 63.8600 67.0560 63.9120 ;
      RECT 0.9000 60.7870 66.1560 63.8600 ;
      RECT 0.0000 60.7390 66.1560 60.7870 ;
      RECT 0.0000 29.0250 66.1560 60.7870 ;
      RECT 0.0000 29.0250 67.0560 60.7390 ;
      RECT 0.9000 29.0250 66.1560 63.8600 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 60.7390 ;
      RECT 0.9000 29.0210 67.0560 29.0250 ;
      RECT 0.9000 27.4250 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.9000 18.3300 66.1560 29.0210 ;
      RECT 0.0000 0.9010 67.0560 9.1560 ;
      RECT 0.9000 9.1560 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 0.9000 0.9010 67.0560 9.1570 ;
      RECT 44.8090 0.9000 67.0560 9.1560 ;
      RECT 44.8090 0.9000 67.0560 9.1560 ;
      RECT 44.8090 0.9000 67.0560 0.9010 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 9.1560 ;
      RECT 46.6670 0.0000 67.0560 0.9000 ;
      RECT 0.0000 72.7280 67.0560 78.3780 ;
      RECT 0.9000 72.6790 67.0560 72.7280 ;
      RECT 0.9000 69.6100 66.1560 72.7280 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 78.4270 66.1560 82.9320 ;
      RECT 0.9000 82.9530 66.1560 86.0970 ;
      RECT 0.9000 78.4270 66.1560 86.0840 ;
  END
END SRAMLP2RW64x8

MACRO SRAMLP2RW64x16
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 88.672 BY 96.013 ;
  SYMMETRY X Y R90 ;

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.7790 0.0000 32.9790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.7790 0.0000 32.9790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.7790 0.0000 32.9790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.7790 0.0000 32.9790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.7790 0.0000 32.9790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[5]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.0960 0.0000 32.2960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.0960 0.0000 32.2960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.0960 0.0000 32.2960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.0960 0.0000 32.2960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.0960 0.0000 32.2960 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[7]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 83.4000 88.6720 83.6000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 83.4000 88.6720 83.6000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 83.4000 88.6720 83.6000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 83.4000 88.6720 83.6000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 83.4000 88.6720 83.6000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 74.5740 88.6720 74.7740 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 74.5740 88.6720 74.7740 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 74.5740 88.6720 74.7740 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 74.5740 88.6720 74.7740 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 74.5740 88.6720 74.7740 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 76.1000 88.6720 76.3000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 76.1000 88.6720 76.3000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 76.1000 88.6720 76.3000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 76.1000 88.6720 76.3000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 76.1000 88.6720 76.3000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 67.3200 88.6720 67.5200 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 67.3200 88.6720 67.5200 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 67.3200 88.6720 67.5200 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 67.3200 88.6720 67.5200 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 67.3200 88.6720 67.5200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 65.7510 88.6720 65.9510 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 65.7510 88.6720 65.9510 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 65.7510 88.6720 65.9510 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 65.7510 88.6720 65.9510 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 65.7510 88.6720 65.9510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.9130 0.0000 21.1130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.9130 0.0000 21.1130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.9130 0.0000 21.1130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.9130 0.0000 21.1130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.9130 0.0000 21.1130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE2

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 32.4990 88.6720 32.6990 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 32.4990 88.6720 32.6990 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 32.4990 88.6720 32.6990 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 32.4990 88.6720 32.6990 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 32.4990 88.6720 32.6990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[5]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 17.2900 88.6720 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 17.2900 88.6720 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 17.2900 88.6720 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 17.2900 88.6720 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 17.2900 88.6720 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 16.8280 88.6720 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 16.8280 88.6720 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 16.8280 88.6720 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 16.8280 88.6720 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 16.8280 88.6720 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 86.8410 95.7130 87.1420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.5410 95.7130 71.8420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.7420 95.7130 16.0430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.5420 95.7130 8.8430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.4420 95.7130 9.7430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9420 95.7130 5.2430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.6430 95.7130 7.9420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.7430 95.7130 7.0420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.6420 95.7130 70.9410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.8410 95.7130 69.1420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.0420 95.7130 13.3430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.3420 95.7130 73.6420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.5430 95.7130 17.8430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.9420 95.7130 68.2420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1430 95.7130 12.4430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.9410 95.7130 86.2420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.5420 95.7130 80.8410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.9410 95.7130 77.2420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.1420 95.7130 21.4430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.0420 95.7130 76.3420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.2430 95.7130 20.5430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.4410 95.7130 81.7420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.6410 95.7130 79.9410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.2420 95.7130 74.5420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4430 95.7130 18.7430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.3420 95.7130 82.6420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.1420 95.7130 75.4410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.3430 95.7130 19.6420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.7420 95.7130 79.0420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.1420 95.7130 66.4420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.3430 95.7130 10.6430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.8420 95.7130 78.1420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.0430 95.7130 22.3430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.7410 95.7130 70.0420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.2410 95.7130 83.5410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2430 95.7130 2.5430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3420 95.7130 1.6420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.6420 95.7130 16.9420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.4410 95.7130 72.7410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8420 95.7130 6.1420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.2430 95.7130 11.5420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.0420 95.7130 67.3410 96.0130 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 18.8920 95.7130 19.1930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.0920 95.7130 71.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.2930 95.7130 15.5930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.8920 95.7130 82.1910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.0930 95.7130 26.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.2920 95.7130 78.5920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.4930 95.7130 22.7930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.9910 95.7130 72.2910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.1920 95.7130 16.4920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.0910 95.7130 80.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.2920 95.7130 24.5930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.4910 95.7130 76.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.6920 95.7130 20.9930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.4910 95.7130 85.7910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.6920 95.7130 29.9920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.3920 95.7130 86.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.5930 95.7130 30.8930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.7910 95.7130 83.0920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.9920 95.7130 27.2930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.5910 95.7130 75.8920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.7920 95.7130 20.0930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.5910 95.7130 66.8920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.7920 95.7130 11.0930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.4910 95.7130 67.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.6920 95.7130 11.9930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.1910 95.7130 70.4910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.3920 95.7130 14.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.8920 95.7130 73.1910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.0930 95.7130 17.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.7910 95.7130 74.0910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.9920 95.7130 18.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.3920 95.7130 68.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.5930 95.7130 12.8930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.8920 95.7130 64.1920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.0930 95.7130 8.3930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.2920 95.7130 33.5930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.3930 95.7130 32.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.8930 95.7130 55.1930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.0920 95.7130 53.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.7920 95.7130 65.0910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.9930 95.7130 9.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.6920 95.7130 38.9930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.1930 95.7130 43.4940 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.4930 95.7130 31.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.4910 95.7130 58.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.6920 95.7130 2.9930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.0910 95.7130 62.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.2920 95.7130 6.5930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.9910 95.7130 63.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.1920 95.7130 7.4930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.8930 95.7130 46.1930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.4920 95.7130 49.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.3930 95.7130 50.6930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.5920 95.7130 48.8920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.7920 95.7130 47.0910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.9920 95.7130 45.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.2920 95.7130 51.5910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.6930 95.7130 47.9940 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.1930 95.7130 52.4940 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.4920 95.7130 40.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.2920 95.7130 42.5910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.0930 95.7130 35.3930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.9930 95.7130 36.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.0920 95.7130 44.3920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.5920 95.7130 39.8920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.8930 95.7130 37.1920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.3930 95.7130 41.6930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.5920 95.7130 57.8910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.7930 95.7130 2.0920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.1910 95.7130 61.4910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.3920 95.7130 5.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.1920 95.7130 34.4930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.2920 95.7130 60.5920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.4930 95.7130 4.7930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.3910 95.7130 59.6910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.5920 95.7130 3.8920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.7920 95.7130 38.0930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.6920 95.7130 56.9920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.7920 95.7130 56.0920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.9920 95.7130 54.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.2920 95.7130 69.5910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.4930 95.7130 13.7920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.9920 95.7130 81.2920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.1930 95.7130 25.4930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.3920 95.7130 77.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.5930 95.7130 21.8930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.5920 95.7130 84.8920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.7930 95.7130 29.0930 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.6910 95.7130 74.9920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.8920 95.7130 28.1920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.6910 95.7130 83.9910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.3920 95.7130 23.6920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.1910 95.7130 79.4910 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.8930 95.7130 10.1920 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.6920 95.7130 65.9910 96.0130 ;
    END
  END VSS

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 86.2600 88.6720 86.4600 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 86.2600 88.6720 86.4600 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 86.2600 88.6720 86.4600 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 86.2600 88.6720 86.4600 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 86.2600 88.6720 86.4600 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS1

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 89.4480 88.6720 89.6480 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 89.4480 88.6720 89.6480 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 89.4480 88.6720 89.6480 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 89.4480 88.6720 89.6480 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 89.4480 88.6720 89.6480 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 86.2720 0.2000 86.4720 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 86.2720 0.2000 86.4720 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 86.2720 0.2000 86.4720 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 86.2720 0.2000 86.4720 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 86.2720 0.2000 86.4720 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 89.4370 0.2000 89.6370 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 89.4370 0.2000 89.6370 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 89.4370 0.2000 89.6370 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 89.4370 0.2000 89.6370 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 89.4370 0.2000 89.6370 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.1770 0.0000 67.3770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.1770 0.0000 67.3770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.1770 0.0000 67.3770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.1770 0.0000 67.3770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.1770 0.0000 67.3770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.9420 95.7130 14.2430 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.8430 95.7130 15.1420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.1420 95.7130 3.4420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.1420 95.7130 84.4410 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.0430 95.7130 4.3420 96.0130 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.0410 95.7130 85.3420 96.0130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.0690 0.0000 55.2690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.0690 0.0000 55.2690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.0690 0.0000 55.2690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.0690 0.0000 55.2690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.0690 0.0000 55.2690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[5]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3860 0.0000 54.5860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.3860 0.0000 54.5860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.3860 0.0000 54.5860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.3860 0.0000 54.5860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.3860 0.0000 54.5860 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[7]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.5940 0.0000 62.7940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.5940 0.0000 62.7940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.5940 0.0000 62.7940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.5940 0.0000 62.7940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.5940 0.0000 62.7940 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[9]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.9090 0.0000 62.1090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.9090 0.0000 62.1090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.9090 0.0000 62.1090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.9090 0.0000 62.1090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.9090 0.0000 62.1090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[9]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.2260 0.0000 61.4260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.2260 0.0000 61.4260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.2260 0.0000 61.4260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.2260 0.0000 61.4260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.2260 0.0000 61.4260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[14]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.5410 0.0000 60.7410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.5410 0.0000 60.7410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.5410 0.0000 60.7410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.5410 0.0000 60.7410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.5410 0.0000 60.7410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[14]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.8580 0.0000 60.0580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.8580 0.0000 60.0580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.8580 0.0000 60.0580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.8580 0.0000 60.0580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.8580 0.0000 60.0580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.1730 0.0000 59.3730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.1730 0.0000 59.3730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.1730 0.0000 59.3730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.1730 0.0000 59.3730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.1730 0.0000 59.3730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[0]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.4900 0.0000 58.6900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.4900 0.0000 58.6900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.4900 0.0000 58.6900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.4900 0.0000 58.6900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.4900 0.0000 58.6900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[13]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4970 0.0000 66.6970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4970 0.0000 66.6970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4970 0.0000 66.6970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4970 0.0000 66.6970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4970 0.0000 66.6970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[3]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.0130 0.0000 66.2130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.0130 0.0000 66.2130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.0130 0.0000 66.2130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.0130 0.0000 66.2130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.0130 0.0000 66.2130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[3]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.3300 0.0000 65.5300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.3300 0.0000 65.5300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.3300 0.0000 65.5300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.3300 0.0000 65.5300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.3300 0.0000 65.5300 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[10]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.6450 0.0000 64.8450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.6450 0.0000 64.8450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.6450 0.0000 64.8450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.6450 0.0000 64.8450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.6450 0.0000 64.8450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[10]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.9620 0.0000 64.1620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.9620 0.0000 64.1620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.9620 0.0000 64.1620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.9620 0.0000 64.1620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.9620 0.0000 64.1620 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.2770 0.0000 63.4770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.2770 0.0000 63.4770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.2770 0.0000 63.4770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.2770 0.0000 63.4770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.2770 0.0000 63.4770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[8]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 9.8200 88.6720 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 9.8200 88.6720 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 9.8200 88.6720 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 9.8200 88.6720 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 9.8200 88.6720 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB2

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4720 85.9200 88.6720 86.1200 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4720 85.9200 88.6720 86.1200 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4720 85.9200 88.6720 86.1200 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4720 85.9200 88.6720 86.1200 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4720 85.9200 88.6720 86.1200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.9360 0.0000 39.1360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.9360 0.0000 39.1360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.9360 0.0000 39.1360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.9360 0.0000 39.1360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.9360 0.0000 39.1360 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[14]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.9140 0.0000 49.1140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.9140 0.0000 49.1140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.9140 0.0000 49.1140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.9140 0.0000 49.1140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.9140 0.0000 49.1140 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[2]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.2290 0.0000 48.4290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.2290 0.0000 48.4290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.2290 0.0000 48.4290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.2290 0.0000 48.4290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.2290 0.0000 48.4290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[2]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.5460 0.0000 47.7460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.5460 0.0000 47.7460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.5460 0.0000 47.7460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.5460 0.0000 47.7460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.5460 0.0000 47.7460 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[15]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.8610 0.0000 47.0610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.8610 0.0000 47.0610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.8610 0.0000 47.0610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.8610 0.0000 47.0610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.8610 0.0000 47.0610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[15]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.1780 0.0000 46.3780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.1780 0.0000 46.3780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.1780 0.0000 46.3780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.1780 0.0000 46.3780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.1780 0.0000 46.3780 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[6]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.4930 0.0000 45.6930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.4930 0.0000 45.6930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.4930 0.0000 45.6930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.4930 0.0000 45.6930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.4930 0.0000 45.6930 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[6]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.8100 0.0000 45.0100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.8100 0.0000 45.0100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.8100 0.0000 45.0100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.8100 0.0000 45.0100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.8100 0.0000 45.0100 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[3]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.7010 0.0000 53.9010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.7010 0.0000 53.9010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.7010 0.0000 53.9010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.7010 0.0000 53.9010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.7010 0.0000 53.9010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[7]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.0180 0.0000 53.2180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.0180 0.0000 53.2180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.0180 0.0000 53.2180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.0180 0.0000 53.2180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.0180 0.0000 53.2180 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.3330 0.0000 52.5330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.3330 0.0000 52.5330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.3330 0.0000 52.5330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.3330 0.0000 52.5330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.3330 0.0000 52.5330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[12]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.6500 0.0000 51.8500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.6500 0.0000 51.8500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.6500 0.0000 51.8500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.6500 0.0000 51.8500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.6500 0.0000 51.8500 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[11]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.9650 0.0000 51.1650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.9650 0.0000 51.1650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.9650 0.0000 51.1650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.9650 0.0000 51.1650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.9650 0.0000 51.1650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[11]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.2820 0.0000 50.4820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.2820 0.0000 50.4820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.2820 0.0000 50.4820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.2820 0.0000 50.4820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.2820 0.0000 50.4820 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.5970 0.0000 49.7970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.5970 0.0000 49.7970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.5970 0.0000 49.7970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.5970 0.0000 49.7970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.5970 0.0000 49.7970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[4]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.8050 0.0000 58.0050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.8050 0.0000 58.0050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.8050 0.0000 58.0050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.8050 0.0000 58.0050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.8050 0.0000 58.0050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[13]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.1220 0.0000 57.3220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.1220 0.0000 57.3220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.1220 0.0000 57.3220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.1220 0.0000 57.3220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.1220 0.0000 57.3220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[1]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.4370 0.0000 56.6370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.4370 0.0000 56.6370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.4370 0.0000 56.6370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.4370 0.0000 56.6370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.4370 0.0000 56.6370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[1]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.7540 0.0000 55.9540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.7540 0.0000 55.9540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.7540 0.0000 55.9540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.7540 0.0000 55.9540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.7540 0.0000 55.9540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O1[5]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.4110 0.0000 31.6110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.4110 0.0000 31.6110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.4110 0.0000 31.6110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.4110 0.0000 31.6110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.4110 0.0000 31.6110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[7]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.7280 0.0000 30.9280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.7280 0.0000 30.9280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.7280 0.0000 30.9280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.7280 0.0000 30.9280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.7280 0.0000 30.9280 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[12]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.0430 0.0000 30.2430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.0430 0.0000 30.2430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.0430 0.0000 30.2430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.0430 0.0000 30.2430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.0430 0.0000 30.2430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[12]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.3600 0.0000 29.5600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.3600 0.0000 29.5600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.3600 0.0000 29.5600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.3600 0.0000 29.5600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.3600 0.0000 29.5600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[11]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.6750 0.0000 28.8750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.6750 0.0000 28.8750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.6750 0.0000 28.8750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.6750 0.0000 28.8750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.6750 0.0000 28.8750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[11]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.2510 0.0000 38.4510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.2510 0.0000 38.4510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.2510 0.0000 38.4510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.2510 0.0000 38.4510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.2510 0.0000 38.4510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[14]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.5680 0.0000 37.7680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.5680 0.0000 37.7680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.5680 0.0000 37.7680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.5680 0.0000 37.7680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.5680 0.0000 37.7680 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[0]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.8830 0.0000 37.0830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.8830 0.0000 37.0830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.8830 0.0000 37.0830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.8830 0.0000 37.0830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.8830 0.0000 37.0830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[0]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.2000 0.0000 36.4000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.2000 0.0000 36.4000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.2000 0.0000 36.4000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.2000 0.0000 36.4000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.2000 0.0000 36.4000 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[13]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.5150 0.0000 35.7150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.5150 0.0000 35.7150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.5150 0.0000 35.7150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.5150 0.0000 35.7150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.5150 0.0000 35.7150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[13]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.8320 0.0000 35.0320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.8320 0.0000 35.0320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.8320 0.0000 35.0320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.8320 0.0000 35.0320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.8320 0.0000 35.0320 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[1]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.1470 0.0000 34.3470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.1470 0.0000 34.3470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.1470 0.0000 34.3470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.1470 0.0000 34.3470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.1470 0.0000 34.3470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[1]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.7230 0.0000 43.9230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.7230 0.0000 43.9230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.7230 0.0000 43.9230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.7230 0.0000 43.9230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.7230 0.0000 43.9230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[3]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.0400 0.0000 43.2400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.0400 0.0000 43.2400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.0400 0.0000 43.2400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.0400 0.0000 43.2400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.0400 0.0000 43.2400 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[10]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.3550 0.0000 42.5550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.3550 0.0000 42.5550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.3550 0.0000 42.5550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.3550 0.0000 42.5550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.3550 0.0000 42.5550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[10]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.6720 0.0000 41.8720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.6720 0.0000 41.8720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.6720 0.0000 41.8720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.6720 0.0000 41.8720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.6720 0.0000 41.8720 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[8]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.9870 0.0000 41.1870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.9870 0.0000 41.1870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.9870 0.0000 41.1870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.9870 0.0000 41.1870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.9870 0.0000 41.1870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[8]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.3040 0.0000 40.5040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.3040 0.0000 40.5040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.3040 0.0000 40.5040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.3040 0.0000 40.5040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.3040 0.0000 40.5040 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[9]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.6190 0.0000 39.8190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.6190 0.0000 39.8190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.6190 0.0000 39.8190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.6190 0.0000 39.8190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.6190 0.0000 39.8190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[9]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB2

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 83.3960 0.2000 83.5960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 83.3960 0.2000 83.5960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 83.3960 0.2000 83.5960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 83.3960 0.2000 83.5960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 74.5780 0.2000 74.7780 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 74.5780 0.2000 74.7780 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 74.5780 0.2000 74.7780 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 74.5780 0.2000 74.7780 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 74.5780 0.2000 74.7780 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 76.0990 0.2000 76.2990 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 76.0990 0.2000 76.2990 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 76.0990 0.2000 76.2990 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 76.0990 0.2000 76.2990 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 76.0990 0.2000 76.2990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 65.7460 0.2000 65.9460 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 65.7460 0.2000 65.9460 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 65.7460 0.2000 65.9460 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 65.7460 0.2000 65.9460 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 65.7460 0.2000 65.9460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[4]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 67.3030 0.2000 67.5030 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 67.3030 0.2000 67.5030 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 67.3030 0.2000 67.5030 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 67.3030 0.2000 67.5030 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 67.3030 0.2000 67.5030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.5000 0.2000 32.7000 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 32.5000 0.2000 32.7000 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 32.5000 0.2000 32.7000 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.5000 0.2000 32.7000 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 32.5000 0.2000 32.7000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[5]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.9920 0.0000 28.1920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.9920 0.0000 28.1920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.9920 0.0000 28.1920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.9920 0.0000 28.1920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.9920 0.0000 28.1920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[4]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.3070 0.0000 27.5070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.3070 0.0000 27.5070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.3070 0.0000 27.5070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.3070 0.0000 27.5070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.3070 0.0000 27.5070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[4]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.6240 0.0000 26.8240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.6240 0.0000 26.8240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.6240 0.0000 26.8240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.6240 0.0000 26.8240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.6240 0.0000 26.8240 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[2]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.9390 0.0000 26.1390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.9390 0.0000 26.1390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.9390 0.0000 26.1390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.9390 0.0000 26.1390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[2]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.2560 0.0000 25.4560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.2560 0.0000 25.4560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.2560 0.0000 25.4560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.2560 0.0000 25.4560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.2560 0.0000 25.4560 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[15]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.5710 0.0010 24.7710 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.5710 0.0010 24.7710 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.5710 0.0000 24.7710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.5710 0.0000 24.7710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.5710 0.0000 24.7710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[15]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.8880 0.0000 24.0880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.8880 0.0000 24.0880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.8880 0.0000 24.0880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.8880 0.0000 24.0880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.8880 0.0000 24.0880 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[6]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.2030 0.0000 23.4030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.2030 0.0000 23.4030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.2030 0.0000 23.4030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.2030 0.0000 23.4030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.2030 0.0000 23.4030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[6]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.4640 0.0000 33.6640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.4640 0.0000 33.6640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.4640 0.0000 33.6640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.4640 0.0000 33.6640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.4640 0.0000 33.6640 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
  END O2[5]
  OBS
    LAYER M1 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 65.1460 87.8720 73.9740 ;
      RECT 0.8000 66.5460 87.8720 66.5510 ;
      RECT 0.8000 33.2990 88.6720 65.1460 ;
      RECT 0.8000 33.2990 88.6720 65.1460 ;
      RECT 0.8000 33.2990 88.6720 65.1460 ;
      RECT 0.8000 33.2990 88.6720 33.3000 ;
      RECT 87.8720 84.2000 88.6720 85.3200 ;
      RECT 21.7130 0.0000 22.6030 0.8000 ;
      RECT 0.0000 87.0720 1.5010 88.8370 ;
      RECT 0.0000 70.9770 87.8720 73.9780 ;
      RECT 0.0000 68.1030 3.0010 68.1200 ;
      RECT 0.0000 90.2370 87.8720 93.2380 ;
      RECT 87.1710 87.0600 88.6720 88.8480 ;
      RECT 87.8720 66.5510 88.6720 66.7200 ;
      RECT 85.6710 65.1460 88.6720 65.1510 ;
      RECT 0.8000 75.4990 88.6720 75.5000 ;
      RECT 0.8000 75.3740 88.6720 75.3780 ;
      RECT 0.8000 73.9780 87.8720 75.3740 ;
      RECT 0.8000 75.5000 87.8720 76.8990 ;
      RECT 0.0000 66.5460 0.8000 66.7030 ;
      RECT 0.0000 75.3780 88.6720 75.4990 ;
      RECT 0.8000 75.3780 87.8720 75.4990 ;
      RECT 0.8000 16.2340 87.8720 18.0900 ;
      RECT 0.0000 16.2280 87.8720 16.2340 ;
      RECT 0.0000 0.0000 20.3130 9.2200 ;
      RECT 0.0000 0.0000 20.3130 0.8000 ;
      RECT 0.0000 10.6210 87.8720 16.2340 ;
      RECT 0.0000 10.6210 87.8720 16.2340 ;
      RECT 0.0000 10.6210 87.8720 16.2340 ;
      RECT 0.0000 10.6210 88.6720 16.2280 ;
      RECT 0.8000 10.6210 87.8720 18.0900 ;
      RECT 0.8000 10.6210 87.8720 18.0900 ;
      RECT 0.8000 10.6210 87.8720 18.0900 ;
      RECT 0.8000 10.6200 88.6720 16.2280 ;
      RECT 0.8000 10.6200 88.6720 16.2280 ;
      RECT 0.8000 10.6200 88.6720 16.2280 ;
      RECT 0.8000 10.6200 88.6720 10.6210 ;
      RECT 0.8000 9.2210 87.8720 10.6200 ;
      RECT 0.0000 31.8990 87.8720 31.9000 ;
      RECT 0.0000 18.1680 87.8720 31.9000 ;
      RECT 0.0000 18.1680 87.8720 31.9000 ;
      RECT 0.0000 18.1680 87.8720 31.9000 ;
      RECT 0.0000 18.1680 88.6720 31.8990 ;
      RECT 0.8000 18.0900 88.6720 31.8990 ;
      RECT 0.8000 18.0900 88.6720 31.8990 ;
      RECT 0.8000 18.0900 88.6720 31.8990 ;
      RECT 0.8000 18.0900 88.6720 18.1680 ;
      RECT 0.8000 31.9000 87.8720 33.2990 ;
      RECT 0.8000 18.1680 87.8720 33.2990 ;
      RECT 0.8000 18.1680 87.8720 33.2990 ;
      RECT 0.8000 18.1680 87.8720 33.2990 ;
      RECT 0.0000 9.2200 87.8720 9.2210 ;
      RECT 0.0000 0.8000 87.8720 9.2210 ;
      RECT 0.0000 0.8000 87.8720 9.2210 ;
      RECT 0.0000 0.8000 87.8720 9.2210 ;
      RECT 0.0000 0.8000 88.6720 9.2200 ;
      RECT 0.8000 0.8000 87.8720 10.6200 ;
      RECT 0.8000 0.8000 87.8720 10.6200 ;
      RECT 0.8000 0.8000 87.8720 10.6200 ;
      RECT 67.9770 0.0000 88.6720 9.2200 ;
      RECT 67.9770 0.0000 88.6720 0.8000 ;
      RECT 0.0000 76.9000 87.8720 85.6720 ;
      RECT 0.0000 76.9000 87.8720 85.6720 ;
      RECT 0.0000 76.9000 87.8720 85.6720 ;
      RECT 0.0000 76.9000 87.8720 85.6720 ;
      RECT 0.0000 76.9000 88.6720 82.8000 ;
      RECT 0.0000 76.8990 87.8720 82.8000 ;
      RECT 0.0000 76.8990 87.8720 76.9000 ;
      RECT 0.8000 75.4990 87.8720 75.5000 ;
      RECT 0.0000 68.1200 88.6720 73.9740 ;
      RECT 0.8000 75.3740 87.8720 75.3780 ;
      RECT 0.0000 90.2480 88.6720 96.0130 ;
      RECT 0.8000 87.0720 87.8720 90.2370 ;
      RECT 0.8000 87.0600 87.8720 90.2370 ;
      RECT 0.8000 87.0600 87.8720 90.2370 ;
      RECT 0.8000 87.0600 87.8720 90.2370 ;
      RECT 0.8000 87.0600 87.8720 90.2370 ;
      RECT 0.8000 87.0600 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 85.6720 87.8720 90.2370 ;
      RECT 0.8000 76.9000 87.8720 87.0600 ;
      RECT 0.8000 76.9000 87.8720 87.0600 ;
      RECT 0.8000 76.9000 87.8720 87.0600 ;
      RECT 0.0000 33.3000 88.6720 65.1460 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
      RECT 0.8000 65.1510 87.8720 73.9740 ;
    LAYER PO ;
      RECT 0.0000 0.0000 88.6720 96.0130 ;
    LAYER M2 ;
      RECT 0.0000 90.3480 88.6720 96.0130 ;
      RECT 0.0000 77.0000 88.6720 82.6960 ;
      RECT 0.0000 76.9990 87.7720 77.0000 ;
      RECT 0.9000 73.8780 87.7720 77.0000 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 87.7720 84.3000 88.6720 85.2200 ;
      RECT 0.0000 84.2960 0.9000 85.5720 ;
      RECT 21.8130 0.0000 22.5030 0.9000 ;
      RECT 0.0000 87.1720 1.5010 88.7370 ;
      RECT 0.0000 90.3370 87.7720 93.3380 ;
      RECT 0.9000 79.6990 88.6720 82.7000 ;
      RECT 87.1710 87.1600 88.6720 88.7480 ;
      RECT 0.0000 68.2200 88.6720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 68.2200 ;
      RECT 0.9000 65.0510 87.7720 73.8740 ;
      RECT 0.9000 65.0510 87.7720 68.2030 ;
      RECT 0.9000 65.0460 88.6720 65.0510 ;
      RECT 0.0000 33.4000 88.6720 65.0460 ;
      RECT 0.9000 33.4000 87.7720 68.2030 ;
      RECT 0.9000 33.4000 88.6720 65.0510 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 33.4000 ;
      RECT 0.9000 31.8000 87.7720 33.3990 ;
      RECT 0.0000 73.8740 87.7720 73.8780 ;
      RECT 0.0000 68.2200 87.7720 73.8780 ;
      RECT 0.9000 73.8780 87.7720 76.9990 ;
      RECT 0.9000 68.2200 87.7720 76.9990 ;
      RECT 0.0000 31.7990 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 88.6720 31.7990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 18.2680 ;
      RECT 0.9000 16.1340 87.7720 18.1900 ;
      RECT 0.0000 16.1280 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 88.6720 16.1280 ;
      RECT 0.9000 10.7210 87.7720 18.1900 ;
      RECT 0.9000 10.7210 87.7720 18.1900 ;
      RECT 0.9000 10.7210 87.7720 18.1900 ;
      RECT 0.0000 0.0000 20.2130 9.1200 ;
      RECT 0.0000 0.0000 20.2130 0.9000 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 10.7210 ;
      RECT 0.9000 9.1210 87.7720 10.7200 ;
      RECT 0.0000 9.1200 87.7720 9.1210 ;
      RECT 0.0000 0.9000 87.7720 9.1210 ;
      RECT 0.0000 0.9000 87.7720 9.1210 ;
      RECT 0.0000 0.9000 87.7720 9.1210 ;
      RECT 0.0000 0.9000 88.6720 9.1200 ;
      RECT 0.9000 0.9000 87.7720 10.7200 ;
      RECT 0.9000 0.9000 87.7720 10.7200 ;
      RECT 0.9000 0.9000 87.7720 10.7200 ;
      RECT 68.0770 0.0000 88.6720 9.1200 ;
      RECT 68.0770 0.0000 88.6720 0.9000 ;
    LAYER M3 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 88.6720 16.1280 ;
      RECT 0.9000 10.7210 87.7720 18.1900 ;
      RECT 0.9000 10.7210 87.7720 18.1900 ;
      RECT 0.9000 10.7210 87.7720 18.1900 ;
      RECT 0.0000 0.0000 20.2130 9.1200 ;
      RECT 0.0000 0.0000 20.2130 0.9000 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 10.7210 ;
      RECT 0.9000 9.1210 87.7720 10.7200 ;
      RECT 0.0000 9.1200 87.7720 9.1210 ;
      RECT 0.0000 0.9000 87.7720 9.1210 ;
      RECT 0.0000 0.9000 87.7720 9.1210 ;
      RECT 0.0000 0.9000 87.7720 9.1210 ;
      RECT 0.0000 0.9000 88.6720 9.1200 ;
      RECT 0.9000 0.9000 87.7720 10.7200 ;
      RECT 0.9000 0.9000 87.7720 10.7200 ;
      RECT 0.9000 0.9000 87.7720 10.7200 ;
      RECT 68.0770 0.0000 88.6720 9.1200 ;
      RECT 68.0770 0.0000 88.6720 0.9000 ;
      RECT 0.0000 90.3480 88.6720 96.0130 ;
      RECT 0.0000 77.0000 88.6720 82.6960 ;
      RECT 0.0000 76.9990 87.7720 77.0000 ;
      RECT 0.9000 73.8780 87.7720 77.0000 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 21.8130 0.0000 22.5030 0.9000 ;
      RECT 0.0000 90.3370 87.7720 93.3380 ;
      RECT 0.0000 87.1720 1.5010 88.7370 ;
      RECT 0.0000 84.2960 0.9000 85.5720 ;
      RECT 0.9000 79.6990 88.6720 82.7000 ;
      RECT 87.1710 87.1600 88.6720 88.7480 ;
      RECT 87.7720 84.3000 88.6720 85.2200 ;
      RECT 0.0000 68.2200 88.6720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 68.2200 ;
      RECT 0.9000 65.0510 87.7720 73.8740 ;
      RECT 0.9000 65.0510 87.7720 68.2030 ;
      RECT 0.9000 65.0460 88.6720 65.0510 ;
      RECT 0.0000 33.4000 88.6720 65.0460 ;
      RECT 0.9000 33.4000 87.7720 68.2030 ;
      RECT 0.9000 33.4000 88.6720 65.0510 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 33.4000 ;
      RECT 0.9000 31.8000 87.7720 33.3990 ;
      RECT 0.0000 73.8740 87.7720 73.8780 ;
      RECT 0.0000 68.2200 87.7720 73.8780 ;
      RECT 0.9000 73.8780 87.7720 76.9990 ;
      RECT 0.9000 68.2200 87.7720 76.9990 ;
      RECT 0.0000 31.7990 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 88.6720 31.7990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 18.2680 ;
      RECT 0.9000 16.1340 87.7720 18.1900 ;
      RECT 0.0000 16.1280 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
    LAYER M4 ;
      RECT 0.9000 65.0460 88.6720 65.0510 ;
      RECT 0.9000 33.4000 88.6720 65.0510 ;
      RECT 0.0000 16.1280 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 88.6720 16.1280 ;
      RECT 0.9000 16.1340 87.7720 18.1900 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 10.7210 ;
      RECT 0.0000 31.7990 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 88.6720 31.7990 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 33.4000 ;
      RECT 0.9000 31.8000 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 10.7210 87.7720 31.7990 ;
      RECT 0.9000 10.7210 87.7720 31.7990 ;
      RECT 0.9000 10.7210 87.7720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 18.2680 ;
      RECT 0.0000 9.1200 87.7720 9.1210 ;
      RECT 0.0000 0.9010 87.7720 9.1210 ;
      RECT 0.0000 0.9010 87.7720 9.1210 ;
      RECT 0.0000 0.9010 87.7720 9.1210 ;
      RECT 0.0000 0.9010 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 0.9010 ;
      RECT 68.0770 0.0000 88.6720 9.1200 ;
      RECT 68.0770 0.0000 88.6720 9.1200 ;
      RECT 68.0770 0.0000 88.6720 0.9000 ;
      RECT 0.0000 90.3480 88.6720 96.0130 ;
      RECT 0.0000 77.0000 88.6720 82.6960 ;
      RECT 0.0000 76.9990 87.7720 77.0000 ;
      RECT 0.9000 73.8780 87.7720 77.0000 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.2200 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 85.5720 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 84.2960 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 88.7370 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 21.8130 0.0000 22.5030 0.9000 ;
      RECT 0.0000 90.3370 87.7720 93.3380 ;
      RECT 0.0000 87.1720 1.5010 88.7370 ;
      RECT 0.0000 84.2960 0.9000 85.5720 ;
      RECT 0.9000 79.6990 88.6720 82.7000 ;
      RECT 87.1710 87.1600 88.6720 88.7480 ;
      RECT 87.7720 84.3000 88.6720 85.2200 ;
      RECT 0.0000 0.0000 20.2130 0.9000 ;
      RECT 0.0000 0.0000 20.2130 9.1200 ;
      RECT 0.0000 0.9000 23.8710 9.1200 ;
      RECT 0.0000 0.9000 23.8710 9.1200 ;
      RECT 0.0000 0.9000 23.8710 9.1200 ;
      RECT 0.0000 0.9000 23.8710 0.9010 ;
      RECT 0.0000 68.2200 88.6720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 68.2200 ;
      RECT 0.0000 73.8740 87.7720 73.8780 ;
      RECT 0.0000 68.2200 87.7720 73.8780 ;
      RECT 0.9000 73.8780 87.7720 76.9990 ;
      RECT 0.9000 68.2200 87.7720 76.9990 ;
      RECT 0.9000 9.1210 87.7720 10.7200 ;
      RECT 0.9000 65.0510 87.7720 73.8740 ;
      RECT 0.9000 65.0510 87.7720 68.2030 ;
      RECT 0.0000 33.4000 88.6720 65.0460 ;
      RECT 0.9000 33.4000 87.7720 68.2030 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 88.6720 96.0130 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 88.6720 96.0130 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 88.6720 96.0130 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 88.6720 96.0130 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 88.6720 96.0130 ;
    LAYER M5 ;
      RECT 0.0000 95.0130 0.6420 96.0130 ;
      RECT 21.8130 0.0000 22.5030 0.9010 ;
      RECT 21.8130 0.0000 22.5030 0.9000 ;
      RECT 21.8130 0.0000 22.5030 0.9010 ;
      RECT 87.8420 95.0130 88.6720 96.0130 ;
      RECT 0.0000 84.2960 0.9000 85.5720 ;
      RECT 0.0000 90.3370 87.7720 93.3380 ;
      RECT 0.0000 87.1720 1.5010 88.7370 ;
      RECT 0.9000 79.6990 88.6720 82.7000 ;
      RECT 87.1710 87.1600 88.6720 88.7480 ;
      RECT 87.7720 84.3000 88.6720 85.2200 ;
      RECT 0.0000 0.9000 23.8710 9.1200 ;
      RECT 0.0000 0.9000 23.8710 9.1200 ;
      RECT 0.0000 0.0000 20.2130 9.1200 ;
      RECT 0.0000 0.9000 23.8710 9.1200 ;
      RECT 0.0000 0.0000 20.2130 9.1200 ;
      RECT 0.0000 0.9000 23.8710 0.9010 ;
      RECT 0.0000 0.0000 20.2130 0.9000 ;
      RECT 0.0000 68.2200 88.6720 73.8740 ;
      RECT 0.0000 73.8740 87.7720 73.8780 ;
      RECT 0.0000 68.2200 87.7720 73.8780 ;
      RECT 0.9000 73.8780 87.7720 76.9990 ;
      RECT 0.9000 68.2200 87.7720 76.9990 ;
      RECT 0.0000 68.2030 87.7720 73.8740 ;
      RECT 0.0000 68.2030 87.7720 68.2200 ;
      RECT 0.9000 65.0510 87.7720 73.8740 ;
      RECT 0.9000 65.0510 87.7720 68.2030 ;
      RECT 0.9000 9.1210 87.7720 10.7200 ;
      RECT 0.0000 16.1280 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 87.7720 16.1340 ;
      RECT 0.0000 10.7210 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 16.1280 ;
      RECT 0.9000 10.7200 88.6720 10.7210 ;
      RECT 0.9000 16.1340 87.7720 18.1900 ;
      RECT 0.0000 31.7990 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 87.7720 31.8000 ;
      RECT 0.0000 18.2680 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 31.7990 ;
      RECT 0.9000 10.7210 87.7720 31.7990 ;
      RECT 0.9000 10.7210 87.7720 31.7990 ;
      RECT 0.9000 10.7210 87.7720 31.7990 ;
      RECT 0.9000 18.1900 88.6720 18.2680 ;
      RECT 0.0000 33.4000 88.6720 65.0460 ;
      RECT 0.9000 33.4000 87.7720 68.2030 ;
      RECT 0.9000 65.0460 88.6720 65.0510 ;
      RECT 0.9000 33.4000 88.6720 65.0510 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 65.0460 ;
      RECT 0.9000 33.3990 88.6720 33.4000 ;
      RECT 0.9000 31.8000 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.9000 18.2680 87.7720 33.3990 ;
      RECT 0.0000 9.1200 87.7720 9.1210 ;
      RECT 0.0000 0.9010 87.7720 9.1210 ;
      RECT 0.0000 0.9010 87.7720 9.1210 ;
      RECT 0.0000 0.9010 87.7720 9.1210 ;
      RECT 0.0000 0.9010 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 9.1200 ;
      RECT 25.4710 0.9000 88.6720 0.9010 ;
      RECT 68.0770 0.0000 88.6720 9.1200 ;
      RECT 68.0770 0.0000 88.6720 9.1200 ;
      RECT 68.0770 0.0000 88.6720 0.9000 ;
      RECT 0.9000 85.2200 87.7720 85.5720 ;
      RECT 0.0000 90.3480 88.6720 95.0130 ;
      RECT 0.0000 77.0000 88.6720 82.6960 ;
      RECT 0.0000 76.9990 87.7720 77.0000 ;
      RECT 0.9000 73.8780 87.7720 77.0000 ;
      RECT 0.9000 87.1720 87.7720 90.3370 ;
      RECT 0.9000 87.1600 87.7720 90.3370 ;
      RECT 0.9000 87.1600 87.7720 90.3370 ;
      RECT 0.9000 87.1600 87.7720 90.3370 ;
      RECT 0.9000 87.1600 87.7720 90.3370 ;
      RECT 0.9000 87.1600 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 85.5720 87.7720 90.3370 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
      RECT 0.9000 82.7000 87.7720 87.1600 ;
  END
END SRAMLP2RW64x16

MACRO SRAMLP2RW64x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 132.461 BY 107.472 ;
  SYMMETRY X Y R90 ;

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 76.0290 0.2000 76.2290 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 76.0290 0.2000 76.2290 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 76.0290 0.2000 76.2290 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 76.0290 0.2000 76.2290 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 76.0290 0.2000 76.2290 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 83.2660 0.2000 83.4660 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 83.2660 0.2000 83.4660 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 83.2660 0.2000 83.4660 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 83.2660 0.2000 83.4660 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 83.2660 0.2000 83.4660 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 92.0790 0.2000 92.2790 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 92.0790 0.2000 92.2790 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 92.0790 0.2000 92.2790 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 92.0790 0.2000 92.2790 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 92.0790 0.2000 92.2790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 84.8670 0.2000 85.0670 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 84.8670 0.2000 85.0670 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 84.8670 0.2000 85.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 84.8670 0.2000 85.0670 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 84.8670 0.2000 85.0670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.9840 0.0000 52.1840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.9840 0.0000 52.1840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.9840 0.0000 52.1840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.9840 0.0000 52.1840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.9840 0.0000 52.1840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[20]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.0880 0.0000 56.2880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.0880 0.0000 56.2880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.0880 0.0000 56.2880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.0880 0.0000 56.2880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.0880 0.0000 56.2880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[18]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7200 0.0000 54.9200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7200 0.0000 54.9200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7200 0.0000 54.9200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7200 0.0000 54.9200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7200 0.0000 54.9200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[7]

  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.7500 0.0020 56.9500 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.7500 0.0020 56.9500 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.7500 0.0020 56.9500 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.7500 0.0020 56.9500 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.7500 0.0020 56.9500 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[18]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.3820 0.0020 55.5820 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.3820 0.0020 55.5820 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.3820 0.0020 55.5820 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.3820 0.0020 55.5820 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.3820 0.0020 55.5820 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.0140 0.0020 54.2140 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.0140 0.0020 54.2140 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.0140 0.0020 54.2140 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.0140 0.0020 54.2140 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.0140 0.0020 54.2140 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[24]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.4560 0.0000 57.6560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.4560 0.0000 57.6560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.4560 0.0000 57.6560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.4560 0.0000 57.6560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.4560 0.0000 57.6560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[17]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.2220 0.0020 62.4220 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.2220 0.0020 62.4220 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.2220 0.0020 62.4220 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.2220 0.0020 62.4220 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.2220 0.0020 62.4220 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.8540 0.0020 61.0540 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.8540 0.0020 61.0540 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.8540 0.0020 61.0540 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.8540 0.0020 61.0540 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.8540 0.0020 61.0540 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.4860 0.0020 59.6860 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.4860 0.0020 59.6860 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.4860 0.0020 59.6860 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.4860 0.0020 59.6860 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.4860 0.0020 59.6860 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 74.4390 132.4610 74.6390 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 74.4390 132.4610 74.6390 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 74.4390 132.4610 74.6390 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 74.4390 132.4610 74.6390 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 74.4390 132.4610 74.6390 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 76.0300 132.4610 76.2300 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 76.0300 132.4610 76.2300 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 76.0300 132.4610 76.2300 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 76.0300 132.4610 76.2300 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 76.0300 132.4610 76.2300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 83.3900 132.4610 83.5900 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 83.3900 132.4610 83.5900 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 83.3900 132.4610 83.5900 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 83.3900 132.4610 83.5900 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 83.3900 132.4610 83.5900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 85.1360 132.4610 85.3360 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 85.1360 132.4610 85.3360 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 85.1360 132.4610 85.3360 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 85.1360 132.4610 85.3360 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 85.1360 132.4610 85.3360 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 92.0780 132.4610 92.2780 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 92.0780 132.4610 92.2780 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 92.0780 132.4610 92.2780 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 92.0780 132.4610 92.2780 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 92.0780 132.4610 92.2780 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.9660 0.0000 21.1660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.9660 0.0000 21.1660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.9660 0.0000 21.1660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.9660 0.0000 21.1660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.9660 0.0000 21.1660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 41.1540 132.4610 41.3540 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 41.1540 132.4610 41.3540 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 41.1540 132.4610 41.3540 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 41.1540 132.4610 41.3540 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 41.1540 132.4610 41.3540 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[5]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 16.9030 132.4610 17.1030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 127.8420 107.1710 128.1410 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.7420 107.1710 129.0420 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.9460 107.1710 1.2460 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.8460 107.1710 2.1450 107.4710 ;
    END
    ANTENNADIFFAREA 10.95167 LAYER M5 ;
    ANTENNADIFFAREA 10.95167 LAYER M6 ;
    ANTENNADIFFAREA 10.95167 LAYER M7 ;
    ANTENNADIFFAREA 10.95167 LAYER M8 ;
    ANTENNADIFFAREA 10.95167 LAYER M9 ;
    ANTENNADIFFAREA 10.95167 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 191.6522 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 191.6522 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.0960 107.1700 4.3970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.1960 107.1700 3.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2970 107.1700 2.5970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.3960 107.1700 1.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9960 107.1700 5.2970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.4960 107.1700 9.7970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.5960 107.1700 8.8970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.6970 107.1700 7.9960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.7970 107.1700 7.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.8970 107.1700 6.1970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.2970 107.1700 11.5960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.3970 107.1700 10.6970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.9960 107.1700 14.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.0970 107.1700 13.3970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.1960 107.1700 12.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.4960 107.1700 18.7970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.5960 107.1700 17.8970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.6960 107.1700 16.9970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.7960 107.1700 16.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.8970 107.1700 15.1960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.1960 107.1700 21.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.2970 107.1700 20.5970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.0960 107.1700 22.3970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.8970 107.1700 24.1960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.9970 107.1700 23.2970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.3970 107.1700 19.6970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.6960 107.1700 25.9960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.5970 107.1700 26.8970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.4960 107.1700 27.7960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.3970 107.1700 28.6970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.7960 107.1700 25.0970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.8970 107.1700 33.1970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.0960 107.1700 31.3970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.2970 107.1700 29.5960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.1970 107.1700 30.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.9960 107.1700 32.2970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.7970 107.1700 34.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.3960 107.1700 37.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.5960 107.1700 35.8970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.4960 107.1700 36.7970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.2960 107.1700 38.5960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.6970 107.1700 34.9960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.7960 107.1700 43.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.1970 107.1700 39.4970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.0960 107.1700 40.3950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.8960 107.1700 42.1960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.9970 107.1700 41.2980 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.2960 107.1700 47.5960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.1970 107.1700 48.4970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.3960 107.1700 46.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.6970 107.1700 43.9970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.4970 107.1700 45.7980 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.5960 107.1700 44.8950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.7960 107.1700 52.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.0960 107.1700 49.3950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.9970 107.1700 50.2980 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.6970 107.1700 52.9970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.8960 107.1700 51.1960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.1960 107.1700 57.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.3960 107.1700 55.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.4960 107.1700 54.7960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.5960 107.1700 53.8960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.2970 107.1700 56.5970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.5950 107.1700 62.8950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.6960 107.1700 61.9960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.7960 107.1700 61.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.9960 107.1700 59.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.0960 107.1700 58.3960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.8970 107.1700 60.1970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.0950 107.1700 67.3950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.1960 107.1700 66.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.2950 107.1700 65.5950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.3950 107.1700 64.6950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.4960 107.1700 63.7960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.5960 107.1700 71.8960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.6970 107.1700 70.9970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.7950 107.1700 70.0950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.8950 107.1700 69.1950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.9960 107.1700 68.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.0950 107.1700 76.3950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.1960 107.1700 75.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.2960 107.1700 74.5960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.3960 107.1700 73.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.9960 107.1700 77.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.4970 107.1700 72.7970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.5960 107.1700 80.8960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.6970 107.1700 79.9970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.7950 107.1700 79.0950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.8950 107.1700 78.1950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.4970 107.1700 81.7970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.8950 107.1700 87.1950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.0950 107.1700 85.3950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.1960 107.1700 84.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.2960 107.1700 83.5960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.3960 107.1700 82.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.9960 107.1700 86.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.3960 107.1700 91.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.4960 107.1700 90.7960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.5960 107.1700 89.8960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.7960 107.1700 88.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.6970 107.1700 88.9970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.9960 107.1700 95.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.0950 107.1700 94.3950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.2950 107.1700 92.5950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.8970 107.1700 96.1970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.1960 107.1700 93.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.2950 107.1700 101.5950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.4950 107.1700 99.7950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.5960 107.1700 98.8960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.6960 107.1700 97.9960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.7960 107.1700 97.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.3960 107.1700 100.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.7970 107.1700 106.0970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.8970 107.1700 105.1970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.9970 107.1700 104.2970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.1970 107.1700 102.4970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.0980 107.1700 103.3980 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.3960 107.1700 109.6960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.4960 107.1700 108.7960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.6960 107.1700 106.9960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.2970 107.1700 110.5970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.5970 107.1700 107.8970 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.6950 107.1700 115.9950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.8950 107.1700 114.1950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.9960 107.1700 113.2960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.0960 107.1700 112.3960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.1960 107.1700 111.4960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.7960 107.1700 115.0960 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.1940 107.1700 120.4940 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.2940 107.1700 119.5940 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.3940 107.1700 118.6940 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.5940 107.1700 116.8940 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.4950 107.1700 117.7950 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.7920 107.1700 124.0920 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.8930 107.1700 123.1930 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.0930 107.1700 121.3930 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.6930 107.1700 124.9930 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.0910 107.1700 130.3910 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.1920 107.1700 129.4920 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.5920 107.1700 125.8920 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.4920 107.1700 126.7920 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.3920 107.1700 127.6920 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.2910 107.1700 128.5910 107.4700 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.9940 107.1700 122.2940 107.4700 ;
    END
    ANTENNADIFFAREA 820.1877 LAYER M5 ;
    ANTENNADIFFAREA 820.1877 LAYER M6 ;
    ANTENNADIFFAREA 820.1877 LAYER M7 ;
    ANTENNADIFFAREA 820.1877 LAYER M8 ;
    ANTENNADIFFAREA 820.1877 LAYER M9 ;
    ANTENNADIFFAREA 820.1877 LAYER MRDL ;
    ANTENNAGATEAREA 32.8836 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 7872.011 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7872.011 LAYER M5 ;
    ANTENNAMAXAREACAR 325.7044 LAYER M5 ;
    ANTENNAGATEAREA 32.8836 LAYER M6 ;
    ANTENNAGATEAREA 32.8836 LAYER M7 ;
    ANTENNAGATEAREA 32.8836 LAYER M8 ;
    ANTENNAGATEAREA 32.8836 LAYER M9 ;
    ANTENNAGATEAREA 32.8836 LAYER MRDL ;
  END VSS

  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.8060 0.0020 46.0060 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.8060 0.0020 46.0060 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.8060 0.0020 46.0060 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.8060 0.0020 46.0060 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.8060 0.0020 46.0060 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[22]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.9100 0.0020 50.1100 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.9100 0.0020 50.1100 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.9100 0.0020 50.1100 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.9100 0.0020 50.1100 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.9100 0.0020 50.1100 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[15]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.6160 0.0000 50.8160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.6160 0.0000 50.8160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.6160 0.0000 50.8160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.6160 0.0000 50.8160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.6160 0.0000 50.8160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[27]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.2480 0.0000 49.4480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.2480 0.0000 49.4480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.2480 0.0000 49.4480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.2480 0.0000 49.4480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.2480 0.0000 49.4480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[15]

  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.6460 0.0020 52.8460 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.6460 0.0020 52.8460 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.6460 0.0020 52.8460 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.6460 0.0020 52.8460 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.6460 0.0020 52.8460 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[20]

  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.2780 0.0020 51.4780 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.2780 0.0020 51.4780 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.2780 0.0020 51.4780 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.2780 0.0020 51.4780 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.2780 0.0020 51.4780 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[27]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.3520 0.0000 53.5520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.3520 0.0000 53.5520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.3520 0.0000 53.5520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.3520 0.0000 53.5520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.3520 0.0000 53.5520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[24]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.4260 0.0000 93.6260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.4260 0.0000 93.6260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.4260 0.0000 93.6260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.4260 0.0000 93.6260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.4260 0.0000 93.6260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[15]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.4640 0.0020 31.6640 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.4640 0.0020 31.6640 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.4640 0.0020 31.6640 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.4640 0.0020 31.6640 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.4640 0.0020 31.6640 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[13]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 96.6200 132.4610 96.8200 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 96.6200 132.4610 96.8200 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 96.6200 132.4610 96.8200 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 96.6200 132.4610 96.8200 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 96.6200 132.4610 96.8200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 97.4500 132.4610 97.6500 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 97.4500 132.4610 97.6500 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 97.4500 132.4610 97.6500 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 97.4500 132.4610 97.6500 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 97.4500 132.4610 97.6500 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS1

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 100.6030 132.4610 100.8030 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 100.6030 132.4610 100.8030 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 100.6030 132.4610 100.8030 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 100.6030 132.4610 100.8030 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 100.6030 132.4610 100.8030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 100.5520 0.2000 100.7520 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 100.5520 0.2000 100.7520 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 100.5520 0.2000 100.7520 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 100.5520 0.2000 100.7520 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 97.4090 0.2000 97.6090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 97.4090 0.2000 97.6090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 97.4090 0.2000 97.6090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 97.4090 0.2000 97.6090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.0060 0.0000 111.2060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.0060 0.0000 111.2060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.0060 0.0000 111.2060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.0060 0.0000 111.2060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.0060 0.0000 111.2060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB2

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 17.3650 132.4610 17.5650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE1

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2610 9.8950 132.4610 10.0950 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB1

  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.8620 0.0020 35.0620 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.8620 0.0020 35.0620 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.8620 0.0020 35.0620 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.8620 0.0020 35.0620 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.8620 0.0020 35.0620 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[28]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.3040 0.0000 38.5040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.3040 0.0000 38.5040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.3040 0.0000 38.5040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.3040 0.0000 38.5040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.3040 0.0000 38.5040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[25]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.9360 0.0000 37.1360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.9360 0.0000 37.1360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.9360 0.0000 37.1360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.9360 0.0000 37.1360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.9360 0.0000 37.1360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[4]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.5680 0.0000 35.7680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.5680 0.0000 35.7680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.5680 0.0000 35.7680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.5680 0.0000 35.7680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.5680 0.0000 35.7680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[11]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.2000 0.0020 34.4000 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.2000 0.0020 34.4000 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.2000 0.0020 34.4000 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.2000 0.0020 34.4000 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.2000 0.0020 34.4000 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[28]

  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.0700 0.0020 43.2700 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.0700 0.0020 43.2700 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.0700 0.0020 43.2700 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.0700 0.0020 43.2700 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.0700 0.0020 43.2700 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[31]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.7020 0.0020 41.9020 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.7020 0.0020 41.9020 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.7020 0.0020 41.9020 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.7020 0.0020 41.9020 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.7020 0.0020 41.9020 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.3340 0.0020 40.5340 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.3340 0.0020 40.5340 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.3340 0.0020 40.5340 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.3340 0.0020 40.5340 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.3340 0.0020 40.5340 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[23]

  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.9660 0.0020 39.1660 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.9660 0.0020 39.1660 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.9660 0.0020 39.1660 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.9660 0.0020 39.1660 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.9660 0.0020 39.1660 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.7760 0.0000 43.9760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.7760 0.0000 43.9760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.7760 0.0000 43.9760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.7760 0.0000 43.9760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.7760 0.0000 43.9760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[26]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.4080 0.0000 42.6080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.4080 0.0000 42.6080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.4080 0.0000 42.6080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.4080 0.0000 42.6080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.4080 0.0000 42.6080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[31]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.0400 0.0000 41.2400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.0400 0.0000 41.2400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.0400 0.0000 41.2400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.0400 0.0000 41.2400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.0400 0.0000 41.2400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[0]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.6720 0.0000 39.8720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.6720 0.0000 39.8720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.6720 0.0000 39.8720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.6720 0.0000 39.8720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.6720 0.0000 39.8720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[23]

  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.4380 0.0020 44.6380 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.4380 0.0020 44.6380 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.4380 0.0020 44.6380 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.4380 0.0020 44.6380 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.4380 0.0020 44.6380 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[26]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.8800 0.0000 48.0800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.8800 0.0000 48.0800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.8800 0.0000 48.0800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.8800 0.0000 48.0800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.8800 0.0000 48.0800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.1440 0.0000 45.3440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.1440 0.0000 45.3440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.1440 0.0000 45.3440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.1440 0.0000 45.3440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.1440 0.0000 45.3440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[22]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.5120 0.0000 46.7120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.5120 0.0000 46.7120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.5120 0.0000 46.7120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.5120 0.0000 46.7120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.5120 0.0000 46.7120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[29]

  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.5420 0.0020 48.7420 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.5420 0.0020 48.7420 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.5420 0.0020 48.7420 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.5420 0.0020 48.7420 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.5420 0.0020 48.7420 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[21]

  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.1750 0.0020 47.3750 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.1750 0.0020 47.3750 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.1750 0.0020 47.3750 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.1750 0.0020 47.3750 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.1750 0.0020 47.3750 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[29]

  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.0220 0.0020 28.2220 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.0220 0.0020 28.2220 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.0220 0.0020 28.2220 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.0220 0.0020 28.2220 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.0220 0.0020 28.2220 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[19]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.6550 0.0020 26.8550 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.6550 0.0020 26.8550 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.6550 0.0020 26.8550 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.6550 0.0020 26.8550 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.6550 0.0020 26.8550 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.2860 0.0020 25.4860 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.2860 0.0020 25.4860 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.2860 0.0020 25.4860 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.2860 0.0020 25.4860 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.2860 0.0020 25.4860 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.3600 0.0020 27.5600 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.3600 0.0020 27.5600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.3600 0.0020 27.5600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.3600 0.0020 27.5600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.3600 0.0020 27.5600 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[19]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.9920 0.0020 26.1920 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.9920 0.0020 26.1920 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.9920 0.0020 26.1920 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.9920 0.0020 26.1920 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.9920 0.0020 26.1920 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[14]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.6240 0.0020 24.8240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.6240 0.0020 24.8240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.6240 0.0020 24.8240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.6240 0.0020 24.8240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.6240 0.0020 24.8240 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[6]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.2560 0.0020 23.4560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.2560 0.0020 23.4560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.2560 0.0020 23.4560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.2560 0.0020 23.4560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.2560 0.0020 23.4560 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[2]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.1260 0.0020 32.3260 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.1260 0.0020 32.3260 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.1260 0.0020 32.3260 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.1260 0.0020 32.3260 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.1260 0.0020 32.3260 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.7580 0.0020 30.9580 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.7580 0.0020 30.9580 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.7580 0.0020 30.9580 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.7580 0.0020 30.9580 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.7580 0.0020 30.9580 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.3900 0.0020 29.5900 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.3900 0.0020 29.5900 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.3900 0.0020 29.5900 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.3900 0.0020 29.5900 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.3900 0.0020 29.5900 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[30]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.8320 0.0020 33.0320 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.8320 0.0020 33.0320 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.8320 0.0020 33.0320 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.8320 0.0020 33.0320 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.8320 0.0020 33.0320 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[1]

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 17.1470 105.9150 17.4460 106.2150 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6470 105.9170 12.9460 106.2170 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.5470 107.1690 4.8460 107.4690 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6460 107.1690 3.9460 107.4690 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6450 107.1710 12.9460 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1450 107.1710 17.4450 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0470 107.1710 18.3470 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7460 107.1710 12.0470 107.4710 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.1420 107.1720 125.4410 107.4720 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.0420 107.1720 126.3410 107.4720 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 191.637 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 191.637 LAYER M5 ;
  END VDDL

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.0960 0.0020 30.2960 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.0960 0.0020 30.2960 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.0960 0.0020 30.2960 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.0960 0.0020 30.2960 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.0960 0.0020 30.2960 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[5]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.7280 0.0020 28.9280 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.7280 0.0020 28.9280 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.7280 0.0020 28.9280 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.7280 0.0020 28.9280 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.7280 0.0020 28.9280 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[30]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.4940 0.0020 33.6940 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.4940 0.0020 33.6940 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.4940 0.0020 33.6940 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.4940 0.0020 33.6940 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.4940 0.0020 33.6940 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.5970 0.0020 37.7970 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.5970 0.0020 37.7970 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.5970 0.0020 37.7970 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.5970 0.0020 37.7970 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.5970 0.0020 37.7970 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.2300 0.0020 36.4300 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.2300 0.0020 36.4300 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.2300 0.0020 36.4300 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.2300 0.0020 36.4300 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.2300 0.0020 36.4300 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[11]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.7640 0.0020 107.9640 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.7640 0.0020 107.9640 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[16]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.1140 0.0000 81.3140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[4]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 103.6600 0.0020 103.8600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.6600 0.0020 103.8600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.6600 0.0020 103.8600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.6600 0.0020 103.8600 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[10]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.5560 0.0020 99.7560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.5560 0.0020 99.7560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.5560 0.0020 99.7560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.5560 0.0020 99.7560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.5560 0.0020 99.7560 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.6340 0.0000 101.8340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.6340 0.0000 101.8340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.6340 0.0000 101.8340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.6340 0.0000 101.8340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.6340 0.0000 101.8340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.2660 0.0000 100.4660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.2660 0.0000 100.4660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.2660 0.0000 100.4660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.2660 0.0000 100.4660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.2660 0.0000 100.4660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[18]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.8980 0.0000 99.0980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.8980 0.0000 99.0980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.8980 0.0000 99.0980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.8980 0.0000 99.0980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.8980 0.0000 99.0980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[7]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.0020 0.0000 103.2020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.0020 0.0000 103.2020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.0020 0.0000 103.2020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.0020 0.0000 103.2020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.0020 0.0000 103.2020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[10]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.3700 0.0000 104.5700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.3700 0.0000 104.5700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.3700 0.0000 104.5700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.3700 0.0000 104.5700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.3700 0.0000 104.5700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[9]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.2920 0.0020 102.4920 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.2920 0.0020 102.4920 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.2920 0.0020 102.4920 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.2920 0.0020 102.4920 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.2920 0.0020 102.4920 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[17]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.3960 0.0020 106.5960 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.3960 0.0020 106.5960 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.3960 0.0020 106.5960 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.3960 0.0020 106.5960 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.3960 0.0020 106.5960 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.0280 0.0020 105.2280 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.0280 0.0020 105.2280 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.0280 0.0020 105.2280 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.0280 0.0020 105.2280 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.0280 0.0020 105.2280 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[9]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.7380 0.0000 105.9380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.7380 0.0000 105.9380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.7380 0.0000 105.9380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.7380 0.0000 105.9380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.7380 0.0000 105.9380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[3]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.5000 0.0020 110.7000 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.5000 0.0020 110.7000 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.5000 0.0020 110.7000 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.5000 0.0020 110.7000 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.5000 0.0020 110.7000 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.1320 0.0020 109.3320 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.1320 0.0020 109.3320 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.1320 0.0020 109.3320 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.1320 0.0020 109.3320 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.1320 0.0020 109.3320 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[8]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.9140 0.0020 24.1140 0.2020 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.6600 0.0020 103.8600 0.2020 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.7640 0.0020 107.9640 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.9140 0.0020 24.1140 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.7640 0.0020 107.9640 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.9140 0.0020 24.1140 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.7640 0.0020 107.9640 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.9140 0.0020 24.1140 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.9140 0.0020 24.1140 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.4740 0.0000 108.6740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.4740 0.0000 108.6740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.4740 0.0000 108.6740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.4740 0.0000 108.6740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.4740 0.0000 108.6740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[8]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.1060 0.0000 107.3060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.1060 0.0000 107.3060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.1060 0.0000 107.3060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.1060 0.0000 107.3060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.1060 0.0000 107.3060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[16]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.8420 0.0000 110.0420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.8420 0.0000 110.0420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.8420 0.0000 110.0420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.8420 0.0000 110.0420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.8420 0.0000 110.0420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.8760 0.0000 86.0760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.8760 0.0000 86.0760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.8760 0.0000 86.0760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.8760 0.0000 86.0760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.8760 0.0000 86.0760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.5080 0.0020 84.7080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.5080 0.0020 84.7080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.5080 0.0020 84.7080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.5080 0.0020 84.7080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.5080 0.0020 84.7080 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277068 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277068 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[23]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.9240 0.0000 88.1240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.9240 0.0000 88.1240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.9240 0.0000 88.1240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.9240 0.0000 88.1240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.9240 0.0000 88.1240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.29115 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29115 LAYER M3 ;
    ANTENNAMAXAREACAR 62.73159 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.94651 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.16094 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.1400 0.0020 83.3400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.1400 0.0020 83.3400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.1400 0.0020 83.3400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.1400 0.0020 83.3400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.1400 0.0020 83.3400 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[25]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.3480 0.0020 91.5480 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.3480 0.0020 91.5480 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.3480 0.0020 91.5480 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.3480 0.0020 91.5480 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.3480 0.0020 91.5480 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[29]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.9800 0.0020 90.1800 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.9800 0.0020 90.1800 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.9800 0.0020 90.1800 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.9800 0.0020 90.1800 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.9800 0.0020 90.1800 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[22]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.6120 0.0020 88.8120 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.6120 0.0020 88.8120 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.6120 0.0020 88.8120 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.6120 0.0020 88.8120 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.6120 0.0020 88.8120 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[26]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6900 0.0000 90.8900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6900 0.0000 90.8900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6900 0.0000 90.8900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6900 0.0000 90.8900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6900 0.0000 90.8900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[29]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.3220 0.0000 89.5220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.3220 0.0000 89.5220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.3220 0.0000 89.5220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.3220 0.0000 89.5220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.3220 0.0000 89.5220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[22]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.0840 0.0020 94.2840 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.0840 0.0020 94.2840 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.0840 0.0020 94.2840 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.0840 0.0020 94.2840 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.0840 0.0020 94.2840 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.7160 0.0020 92.9160 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.7160 0.0020 92.9160 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.7160 0.0020 92.9160 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.7160 0.0020 92.9160 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.7160 0.0020 92.9160 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[21]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.7940 0.0000 94.9940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.7940 0.0000 94.9940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.7940 0.0000 94.9940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.7940 0.0000 94.9940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.7940 0.0000 94.9940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[27]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.0580 0.0000 92.2580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.0580 0.0000 92.2580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.0580 0.0000 92.2580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.0580 0.0000 92.2580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.0580 0.0000 92.2580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[21]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.1620 0.0000 96.3620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.1620 0.0000 96.3620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.1620 0.0000 96.3620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.1620 0.0000 96.3620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.1620 0.0000 96.3620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[20]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.1890 0.0020 98.3890 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.1890 0.0020 98.3890 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.1890 0.0020 98.3890 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.1890 0.0020 98.3890 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.1890 0.0020 98.3890 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277668 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277668 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[24]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.8200 0.0020 97.0200 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.8200 0.0020 97.0200 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.8200 0.0020 97.0200 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.8200 0.0020 97.0200 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.8200 0.0020 97.0200 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[20]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.5300 0.0000 97.7300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.5300 0.0000 97.7300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.5300 0.0000 97.7300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.5300 0.0000 97.7300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.5300 0.0000 97.7300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[24]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.4520 0.0020 95.6520 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.4520 0.0020 95.6520 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.4520 0.0020 95.6520 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.4520 0.0020 95.6520 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.4520 0.0020 95.6520 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277068 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277068 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[27]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.9240 0.0020 101.1240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.9240 0.0020 101.1240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.9240 0.0020 101.1240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.9240 0.0020 101.1240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.9240 0.0020 101.1240 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[18]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.5380 0.0000 71.7380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.5380 0.0000 71.7380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.5380 0.0000 71.7380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.5380 0.0000 71.7380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.5380 0.0000 71.7380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[19]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.3000 0.0020 76.5000 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.3000 0.0020 76.5000 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.3000 0.0020 76.5000 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.3000 0.0020 76.5000 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.3000 0.0020 76.5000 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.6420 0.0000 75.8420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.6420 0.0000 75.8420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.6420 0.0000 75.8420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.6420 0.0000 75.8420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.6420 0.0000 75.8420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.9320 0.0020 75.1320 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.9320 0.0020 75.1320 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.9320 0.0020 75.1320 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.9320 0.0020 75.1320 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.9320 0.0020 75.1320 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.6680 0.0020 77.8680 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.6680 0.0020 77.8680 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.6680 0.0020 77.8680 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.6680 0.0020 77.8680 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.6680 0.0020 77.8680 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.0100 0.0000 77.2100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.0100 0.0000 77.2100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.0100 0.0000 77.2100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.0100 0.0000 77.2100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.0100 0.0000 77.2100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.7720 0.0020 81.9720 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.7720 0.0020 81.9720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.7720 0.0020 81.9720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.7720 0.0020 81.9720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.7720 0.0020 81.9720 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.4040 0.0020 80.6040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.4040 0.0020 80.6040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.4040 0.0020 80.6040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.4040 0.0020 80.6040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.4040 0.0020 80.6040 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.0360 0.0020 79.2360 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.0360 0.0020 79.2360 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.0360 0.0020 79.2360 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.0360 0.0020 79.2360 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.0360 0.0020 79.2360 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[28]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.1700 0.0000 70.3700 0.2000 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.1140 0.0000 81.3140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.1700 0.0000 70.3700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.1140 0.0000 81.3140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.1700 0.0000 70.3700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.1140 0.0000 81.3140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.1700 0.0000 70.3700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.1700 0.0000 70.3700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.1140 0.0000 81.3140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.7460 0.0000 79.9460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.7460 0.0000 79.9460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.7460 0.0000 79.9460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.7460 0.0000 79.9460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.7460 0.0000 79.9460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.3780 0.0000 78.5780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.3780 0.0000 78.5780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.3780 0.0000 78.5780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.3780 0.0000 78.5780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.3780 0.0000 78.5780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[28]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.4820 0.0000 82.6820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.4820 0.0000 82.6820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.4820 0.0000 82.6820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.4820 0.0000 82.6820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.4820 0.0000 82.6820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[25]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.5860 0.0000 86.7860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.5860 0.0000 86.7860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.5860 0.0000 86.7860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.5860 0.0000 86.7860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.5860 0.0000 86.7860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[31]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.2180 0.0000 85.4180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.2180 0.0000 85.4180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.2180 0.0000 85.4180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.2180 0.0000 85.4180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.2180 0.0000 85.4180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.8500 0.0000 84.0500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.8500 0.0000 84.0500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.8500 0.0000 84.0500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.8500 0.0000 84.0500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.8500 0.0000 84.0500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[23]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.2440 0.0020 87.4440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.2440 0.0020 87.4440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.2440 0.0020 87.4440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.2440 0.0020 87.4440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.2440 0.0020 87.4440 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[31]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.5600 0.0000 61.7600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.5600 0.0000 61.7600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.5600 0.0000 61.7600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.5600 0.0000 61.7600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.5600 0.0000 61.7600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.1920 0.0000 60.3920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.1920 0.0000 60.3920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.1920 0.0000 60.3920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.1920 0.0000 60.3920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.1920 0.0000 60.3920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.8240 0.0000 59.0240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.8240 0.0000 59.0240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.8240 0.0000 59.0240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.8240 0.0000 59.0240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.8240 0.0000 59.0240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.1180 0.0020 58.3180 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.1180 0.0020 58.3180 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.1180 0.0020 58.3180 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.1180 0.0020 58.3180 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.1180 0.0020 58.3180 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[17]

  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.5900 0.0020 63.7900 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.5900 0.0020 63.7900 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.5900 0.0020 63.7900 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.5900 0.0020 63.7900 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.5900 0.0020 63.7900 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[16]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.9280 0.0000 63.1280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.9280 0.0000 63.1280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.9280 0.0000 63.1280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.9280 0.0000 63.1280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.9280 0.0000 63.1280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[16]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.3210 0.0020 66.5210 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.3210 0.0020 66.5210 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.3210 0.0020 66.5210 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.3210 0.0020 66.5210 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.3210 0.0020 66.5210 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.9580 0.0020 65.1580 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.9580 0.0020 65.1580 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.9580 0.0020 65.1580 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.9580 0.0020 65.1580 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.9580 0.0020 65.1580 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.6640 0.0000 65.8640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.6640 0.0000 65.8640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.6640 0.0000 65.8640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.6640 0.0000 65.8640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6640 0.0000 65.8640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.2960 0.0000 64.4960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.2960 0.0000 64.4960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.2960 0.0000 64.4960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.2960 0.0000 64.4960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.2960 0.0000 64.4960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.4600 0.0020 69.6600 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.4600 0.0020 69.6600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.4600 0.0020 69.6600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.4600 0.0020 69.6600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.4600 0.0020 69.6600 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.0920 0.0020 68.2920 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.0920 0.0020 68.2920 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.0920 0.0020 68.2920 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.0920 0.0020 68.2920 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.0920 0.0020 68.2920 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.4340 0.0000 67.6340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.4340 0.0000 67.6340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.4340 0.0000 67.6340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.4340 0.0000 67.6340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.4340 0.0000 67.6340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8020 0.0000 69.0020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8020 0.0000 69.0020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8020 0.0000 69.0020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8020 0.0000 69.0020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8020 0.0000 69.0020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.8280 0.0020 71.0280 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.8280 0.0020 71.0280 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.8280 0.0020 71.0280 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.8280 0.0020 71.0280 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.8280 0.0020 71.0280 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[14]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.5640 0.0020 73.7640 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.5640 0.0020 73.7640 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.5640 0.0020 73.7640 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.5640 0.0020 73.7640 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.5640 0.0020 73.7640 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[30]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.1960 0.0020 72.3960 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.1960 0.0020 72.3960 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.1960 0.0020 72.3960 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.1960 0.0020 72.3960 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.1960 0.0020 72.3960 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[19]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.2740 0.0000 74.4740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.2740 0.0000 74.4740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.2740 0.0000 74.4740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.2740 0.0000 74.4740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.2740 0.0000 74.4740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.9060 0.0000 73.1060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.9060 0.0000 73.1060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.9060 0.0000 73.1060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.9060 0.0000 73.1060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.9060 0.0000 73.1060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[30]

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.43012 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43012 LAYER M4 ;
    ANTENNAMAXAREACAR 13.71244 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.85361 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.33244 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.33244 LAYER M4 ;
    ANTENNAMAXAREACAR 13.19736 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.62924 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE2

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 41.2200 0.2000 41.4200 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 41.2200 0.2000 41.4200 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 41.2200 0.2000 41.4200 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 41.2200 0.2000 41.4200 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 41.2200 0.2000 41.4200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.021 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.99267 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.99267 LAYER M1 ;
    ANTENNAGATEAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAMAXAREACAR 54.48593 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 61.70138 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 68.91637 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.13087 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[5]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 74.4390 0.2000 74.6390 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 74.4390 0.2000 74.6390 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 74.4390 0.2000 74.6390 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 74.4390 0.2000 74.6390 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 74.4390 0.2000 74.6390 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.2527 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2527 LAYER M3 ;
    ANTENNAMAXAREACAR 26.83681 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 30.97712 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 35.11715 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[4]
  OBS
    LAYER M2 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 91.3790 131.5610 99.8520 ;
      RECT 0.9000 91.3790 131.5610 99.8520 ;
      RECT 0.9000 86.0360 131.5610 99.8520 ;
      RECT 0.9000 86.0360 131.5610 99.8520 ;
      RECT 67.2210 0.9000 67.3920 0.9020 ;
      RECT 0.0000 101.4520 131.5610 104.4530 ;
      RECT 0.0000 92.9790 3.0010 96.7090 ;
      RECT 0.0000 91.3780 3.0010 91.3790 ;
      RECT 0.0000 98.3090 1.5010 99.8520 ;
      RECT 0.9000 79.6890 132.4610 82.6900 ;
      RECT 21.8660 0.0000 22.5560 0.9000 ;
      RECT 67.2210 0.9000 67.3920 1.0510 ;
      RECT 85.4080 0.9000 86.5440 1.2010 ;
      RECT 130.9600 92.9790 132.4610 95.9200 ;
      RECT 130.9600 98.3500 132.4610 99.9030 ;
      RECT 131.5610 84.2900 132.4610 84.4360 ;
      RECT 131.5610 92.9780 132.4610 92.9790 ;
      RECT 0.0000 0.0000 20.2660 0.9000 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 0.9020 ;
      RECT 0.0000 40.4540 131.5610 40.5200 ;
      RECT 0.9000 42.0540 132.4610 42.1200 ;
      RECT 0.9000 40.5200 131.5610 42.0540 ;
      RECT 0.0000 42.1200 132.4610 73.7390 ;
      RECT 0.9000 73.7390 131.5610 76.9290 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 132.4610 40.4540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 0.9020 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 0.9000 ;
      RECT 0.0000 86.0360 132.4610 91.3780 ;
      RECT 0.0000 85.7670 131.5610 86.0360 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.0000 101.5030 132.4610 107.4720 ;
      RECT 0.0000 76.9300 132.4610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 76.9300 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 73.7390 131.5610 82.5660 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
    LAYER M1 ;
      RECT 67.1210 0.8000 67.4920 0.8020 ;
      RECT 0.0000 76.8290 3.0010 76.8300 ;
      RECT 0.0000 93.8080 131.6610 96.8090 ;
      RECT 0.0000 84.0660 0.8000 84.2670 ;
      RECT 0.0000 98.2090 1.5010 99.9520 ;
      RECT 0.0000 75.2390 0.8000 75.4290 ;
      RECT 0.0000 101.3520 131.6610 104.3530 ;
      RECT 21.7660 0.0000 22.6560 0.8000 ;
      RECT 67.1210 0.8000 67.4920 1.1010 ;
      RECT 85.3080 0.8000 86.6440 1.1010 ;
      RECT 129.4600 82.6660 132.4610 82.7900 ;
      RECT 130.9600 98.2500 132.4610 100.0030 ;
      RECT 131.6610 84.1900 132.4610 84.5360 ;
      RECT 131.6610 75.2390 132.4610 75.4300 ;
      RECT 0.0000 0.0000 20.3660 9.2950 ;
      RECT 0.0000 0.0000 20.3660 9.2950 ;
      RECT 0.0000 0.8000 22.6560 9.2950 ;
      RECT 0.0000 0.8000 22.6560 9.2950 ;
      RECT 0.0000 0.8000 22.6560 0.8020 ;
      RECT 0.0000 0.0000 20.3660 0.8000 ;
      RECT 0.0000 85.9360 132.4610 91.4780 ;
      RECT 0.0000 85.6670 131.6610 91.4780 ;
      RECT 0.0000 85.6670 131.6610 91.4780 ;
      RECT 0.0000 85.6670 131.6610 91.4780 ;
      RECT 0.0000 85.6670 131.6610 85.9360 ;
      RECT 0.0000 91.4780 131.6610 91.4790 ;
      RECT 0.0000 85.9360 131.6610 91.4790 ;
      RECT 0.0000 85.9360 131.6610 91.4790 ;
      RECT 0.0000 85.9360 131.6610 91.4790 ;
      RECT 0.8000 91.4790 131.6610 92.8780 ;
      RECT 0.0000 16.3030 131.6610 16.3090 ;
      RECT 0.0000 10.6960 131.6610 16.3090 ;
      RECT 0.0000 10.6960 131.6610 16.3090 ;
      RECT 0.0000 10.6960 131.6610 16.3090 ;
      RECT 0.0000 10.6960 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 16.3030 ;
      RECT 0.8000 10.6950 132.4610 10.6960 ;
      RECT 0.8000 9.2960 131.6610 10.6950 ;
      RECT 0.0000 42.0200 132.4610 73.8390 ;
      RECT 0.8000 41.9540 132.4610 73.8390 ;
      RECT 0.8000 41.9540 132.4610 73.8390 ;
      RECT 0.8000 41.9540 132.4610 73.8390 ;
      RECT 0.8000 41.9540 132.4610 42.0200 ;
      RECT 0.8000 40.6200 131.6610 41.9540 ;
      RECT 0.0000 40.5540 131.6610 40.6200 ;
      RECT 0.0000 18.2430 131.6610 40.6200 ;
      RECT 0.0000 18.2430 131.6610 40.6200 ;
      RECT 0.0000 18.2430 131.6610 40.6200 ;
      RECT 0.0000 18.2430 132.4610 40.5540 ;
      RECT 0.8000 18.2430 131.6610 41.9540 ;
      RECT 0.8000 18.2430 131.6610 41.9540 ;
      RECT 0.8000 18.2430 131.6610 41.9540 ;
      RECT 0.8000 18.1650 132.4610 40.5540 ;
      RECT 0.8000 18.1650 132.4610 40.5540 ;
      RECT 0.8000 18.1650 132.4610 40.5540 ;
      RECT 0.8000 18.1650 132.4610 18.2430 ;
      RECT 0.8000 16.3090 131.6610 18.1650 ;
      RECT 0.0000 9.2950 131.6610 9.2960 ;
      RECT 0.0000 0.8020 131.6610 9.2960 ;
      RECT 0.0000 0.8020 131.6610 9.2960 ;
      RECT 0.0000 0.8020 131.6610 9.2960 ;
      RECT 0.0000 0.8020 132.4610 9.2950 ;
      RECT 111.3000 0.8000 132.4610 9.2950 ;
      RECT 111.3000 0.8000 132.4610 9.2950 ;
      RECT 111.3000 0.8000 132.4610 0.8020 ;
      RECT 111.8060 0.0000 132.4610 9.2950 ;
      RECT 111.8060 0.0000 132.4610 9.2950 ;
      RECT 111.8060 0.0000 132.4610 0.8000 ;
      RECT 0.0000 92.8790 132.4610 96.0200 ;
      RECT 0.8000 92.8780 132.4610 92.8790 ;
      RECT 0.0000 76.8300 132.4610 82.6660 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 82.6660 131.6610 85.6670 ;
      RECT 0.8000 84.0660 131.6610 84.1900 ;
      RECT 0.0000 101.4030 132.4610 107.4720 ;
      RECT 0.8000 98.2090 131.6610 101.3520 ;
      RECT 0.8000 98.2090 131.6610 101.3520 ;
      RECT 0.8000 98.2090 131.6610 101.3520 ;
      RECT 0.8000 98.2500 131.6610 101.3520 ;
      RECT 0.8000 98.2090 131.6610 101.3520 ;
      RECT 0.8000 98.2090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 96.8090 131.6610 101.3520 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
      RECT 0.8000 73.8390 131.6610 82.6660 ;
    LAYER PO ;
      RECT 0.0000 0.0000 132.4610 107.4720 ;
    LAYER M3 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 132.4610 40.4540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 0.9020 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 0.9000 ;
      RECT 0.0000 86.0360 132.4610 91.3780 ;
      RECT 0.0000 85.7670 131.5610 86.0360 ;
      RECT 0.0000 101.5030 132.4610 107.4720 ;
      RECT 0.0000 98.3500 131.5610 99.9030 ;
      RECT 0.0000 92.9790 131.5610 101.5030 ;
      RECT 0.0000 95.9200 131.5610 99.9030 ;
      RECT 0.0000 92.9790 131.5610 99.9030 ;
      RECT 0.0000 95.9200 131.5610 99.9030 ;
      RECT 0.0000 92.9790 131.5610 99.9030 ;
      RECT 0.0000 92.9790 131.5610 99.9030 ;
      RECT 0.0000 95.9200 131.5610 99.9030 ;
      RECT 0.0000 95.9200 131.5610 99.9030 ;
      RECT 0.0000 95.9200 131.5610 99.9030 ;
      RECT 0.9000 91.3790 131.5610 98.3500 ;
      RECT 0.9000 86.0360 131.5610 98.3500 ;
      RECT 0.9000 86.0360 131.5610 98.3500 ;
      RECT 0.9000 86.0360 131.5610 98.3500 ;
      RECT 0.9000 86.0360 131.5610 95.9200 ;
      RECT 0.0000 76.9300 132.4610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 76.9300 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 73.7390 131.5610 82.5660 ;
      RECT 67.2210 0.9000 67.3920 0.9020 ;
      RECT 21.8660 0.0000 22.5560 0.9000 ;
      RECT 85.4080 0.9000 86.5440 0.9020 ;
      RECT 0.0000 91.3780 3.0010 91.3790 ;
      RECT 0.9000 79.6890 132.4610 82.6900 ;
      RECT 67.2210 0.9000 67.3920 1.0510 ;
      RECT 85.4080 0.9000 86.5440 1.2010 ;
      RECT 130.9600 98.3500 132.4610 99.9030 ;
      RECT 130.9600 92.9780 132.4610 95.9200 ;
      RECT 131.5610 84.2900 132.4610 84.4360 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 0.9020 ;
      RECT 0.0000 0.0000 20.2660 0.9000 ;
      RECT 0.9000 73.7390 131.5610 76.9290 ;
      RECT 0.0000 40.4540 131.5610 40.5200 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 42.1200 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 42.1200 ;
      RECT 0.9000 40.5200 131.5610 42.0540 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
    LAYER M4 ;
      RECT 0.9000 79.6890 132.4610 82.6900 ;
      RECT 67.2210 0.9000 67.3920 1.0510 ;
      RECT 85.4080 0.9000 86.5440 1.2010 ;
      RECT 130.9600 92.9790 132.4610 95.9200 ;
      RECT 130.9600 98.3500 132.4610 99.9030 ;
      RECT 131.5610 84.2900 132.4610 84.4360 ;
      RECT 131.5610 92.9780 132.4610 92.9790 ;
      RECT 0.0000 0.0000 20.2660 0.9000 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 0.9020 ;
      RECT 0.0000 40.4540 131.5610 40.5200 ;
      RECT 0.9000 42.0540 132.4610 42.1200 ;
      RECT 0.9000 40.5200 131.5610 42.0540 ;
      RECT 0.0000 42.1200 132.4610 73.7390 ;
      RECT 0.9000 73.7390 131.5610 76.9290 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 132.4610 40.4540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 0.9020 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 0.9000 ;
      RECT 0.0000 86.0360 132.4610 91.3780 ;
      RECT 0.0000 85.7670 131.5610 86.0360 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.9000 86.0360 131.5610 92.9790 ;
      RECT 0.0000 101.5030 132.4610 107.4720 ;
      RECT 0.0000 76.9300 132.4610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 76.9300 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 73.7390 131.5610 82.5660 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 98.3500 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 96.7090 131.5610 101.4520 ;
      RECT 0.9000 91.3790 131.5610 99.8520 ;
      RECT 0.9000 91.3790 131.5610 99.8520 ;
      RECT 0.9000 86.0360 131.5610 99.8520 ;
      RECT 0.9000 86.0360 131.5610 99.8520 ;
      RECT 67.2210 0.9000 67.3920 0.9020 ;
      RECT 21.8660 0.0000 22.5560 0.9000 ;
      RECT 85.4080 0.9000 86.5440 0.9020 ;
      RECT 0.0000 101.4520 131.5610 104.4530 ;
      RECT 0.0000 92.9790 3.0010 96.7090 ;
      RECT 0.0000 91.3780 3.0010 91.3790 ;
      RECT 0.0000 98.3090 1.5010 99.8520 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 132.4610 107.4720 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 132.4610 107.4720 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 132.4610 107.4720 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 132.4610 107.4720 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 132.4610 107.4720 ;
    LAYER M5 ;
      RECT 0.0000 106.4710 0.2460 107.4720 ;
      RECT 0.0000 106.4700 0.2460 107.4720 ;
      RECT 0.0000 106.4700 0.2460 107.4720 ;
      RECT 0.0000 106.4700 0.2460 107.4720 ;
      RECT 67.2210 0.9000 67.3920 0.9020 ;
      RECT 0.0000 105.2170 2.9460 106.4700 ;
      RECT 0.0000 106.4700 0.6960 106.4710 ;
      RECT 0.0000 105.2170 2.9460 106.4700 ;
      RECT 0.0000 105.2170 0.6960 106.4710 ;
      RECT 0.0000 105.2170 2.9460 106.4700 ;
      RECT 0.0000 105.2170 0.6960 106.4710 ;
      RECT 0.0000 105.2170 2.9460 106.4700 ;
      RECT 21.8660 0.0000 22.5560 0.9000 ;
      RECT 85.4080 0.9000 86.5440 0.9020 ;
      RECT 131.0910 106.4700 132.4610 107.4720 ;
      RECT 0.0000 106.4690 2.9460 106.4700 ;
      RECT 13.6460 105.2170 16.4470 106.4700 ;
      RECT 0.0000 98.3500 1.5010 99.8520 ;
      RECT 0.0000 98.3090 0.9000 98.3500 ;
      RECT 0.9000 91.3790 131.5610 92.9780 ;
      RECT 13.6460 104.9690 16.4470 106.4700 ;
      RECT 67.2210 0.9000 67.3920 1.0510 ;
      RECT 85.4080 0.9000 86.5440 1.2010 ;
      RECT 130.9600 92.9790 132.4610 95.9200 ;
      RECT 130.9600 98.3500 132.4610 99.8520 ;
      RECT 131.5610 92.9780 132.4610 92.9790 ;
      RECT 131.5610 84.2900 132.4610 84.4360 ;
      RECT 131.5610 99.8520 132.4610 99.9030 ;
      RECT 0.0000 0.0000 20.2660 0.9000 ;
      RECT 0.0000 105.2150 16.4470 105.2170 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.0000 20.2660 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 9.1950 ;
      RECT 0.0000 0.9000 22.5560 0.9020 ;
      RECT 0.0000 10.7960 132.4610 16.2030 ;
      RECT 0.0000 16.2030 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.0000 10.7960 131.5610 16.2090 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 16.2030 ;
      RECT 0.9000 10.7950 132.4610 10.7960 ;
      RECT 0.9000 9.1960 131.5610 10.7950 ;
      RECT 0.9000 16.2090 131.5610 18.2650 ;
      RECT 0.0000 85.7670 131.5610 86.0360 ;
      RECT 0.0000 76.9290 131.5610 76.9300 ;
      RECT 0.0000 101.5030 16.4470 105.2170 ;
      RECT 0.0000 40.4540 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 131.5610 40.5200 ;
      RECT 0.0000 18.3430 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 40.4540 ;
      RECT 0.9000 18.2650 132.4610 18.3430 ;
      RECT 0.0000 42.1200 132.4610 73.7390 ;
      RECT 0.9000 73.7390 131.5610 76.9290 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 73.7390 ;
      RECT 0.9000 42.0540 132.4610 42.1200 ;
      RECT 0.9000 40.5200 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.9000 18.3430 131.5610 42.0540 ;
      RECT 0.0000 95.9200 131.5610 96.7090 ;
      RECT 0.0000 92.9790 131.5610 96.7090 ;
      RECT 0.0000 92.9790 131.5610 96.7090 ;
      RECT 0.0000 92.9790 131.5610 96.7090 ;
      RECT 0.0000 92.9790 131.5610 96.7090 ;
      RECT 0.0000 92.9790 131.5610 95.9200 ;
      RECT 0.9000 98.3500 131.5610 99.8520 ;
      RECT 0.9000 96.7090 131.5610 99.8520 ;
      RECT 0.9000 96.7090 131.5610 99.8520 ;
      RECT 0.9000 95.9200 131.5610 99.8520 ;
      RECT 0.9000 95.9200 131.5610 99.8520 ;
      RECT 0.9000 95.9200 131.5610 99.8520 ;
      RECT 0.9000 95.9200 131.5610 99.8520 ;
      RECT 0.9000 95.9200 131.5610 99.8520 ;
      RECT 0.9000 98.3090 131.5610 98.3500 ;
      RECT 0.0000 105.2170 11.9470 106.4690 ;
      RECT 5.5460 106.4690 11.9470 106.4700 ;
      RECT 0.0000 101.4520 131.5610 101.5030 ;
      RECT 0.9000 98.3500 131.5610 101.5030 ;
      RECT 0.0000 101.5030 132.4610 105.2150 ;
      RECT 18.1460 105.2150 132.4610 106.4700 ;
      RECT 18.1460 101.5030 132.4610 106.4700 ;
      RECT 18.1460 101.5030 132.4610 106.4700 ;
      RECT 0.0000 9.1950 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 131.5610 9.1960 ;
      RECT 0.0000 0.9020 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 9.1950 ;
      RECT 111.4000 0.9000 132.4610 0.9020 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 9.1950 ;
      RECT 111.9060 0.0000 132.4610 0.9000 ;
      RECT 0.0000 76.9300 132.4610 82.5660 ;
      RECT 0.0000 76.9290 131.5610 82.5660 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 86.0360 ;
      RECT 0.9000 82.6900 131.5610 85.7670 ;
      RECT 0.9000 84.2900 131.5610 84.4360 ;
      RECT 0.9000 82.5660 132.4610 82.6900 ;
      RECT 0.9000 73.7390 131.5610 82.5660 ;
      RECT 0.0000 91.3780 131.5610 91.3790 ;
      RECT 0.0000 86.0360 132.4610 91.3780 ;
      RECT 0.9000 92.9780 131.5610 92.9790 ;
  END
END SRAMLP2RW64x32

MACRO SRAMLP2RW128x4
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 54.606 BY 139.784 ;
  SYMMETRY X Y R90 ;

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0000 17.1170 0.2000 17.3170 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0000 16.7390 0.2000 16.9390 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB2

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 129.3710 0.2000 129.5710 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 129.3710 0.2000 129.5710 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 129.3710 0.2000 129.5710 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 129.3710 0.2000 129.5710 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS2

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 110.4680 54.6060 110.6680 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 110.4680 54.6060 110.6680 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 110.4680 54.6060 110.6680 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 110.4680 54.6060 110.6680 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 110.4680 54.6060 110.6680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[3]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.4240 0.0000 25.6240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.7920 0.0000 26.9920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[1]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.4740 0.0000 27.6740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.4740 0.0000 27.6740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.4740 0.0000 27.6740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.4740 0.0000 27.6740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.4740 0.0000 27.6740 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.268488 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.268488 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.5620 0.0000 28.7620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.5620 0.0000 28.7620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.5620 0.0000 28.7620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.5620 0.0000 28.7620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.5620 0.0000 28.7620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[3]

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.4000 0.0000 20.6000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.4000 0.0000 20.6000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.4000 0.0000 20.6000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.4000 0.0000 20.6000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.4000 0.0000 20.6000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB2

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.9300 0.0000 30.1300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.9300 0.0000 30.1300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.9300 0.0000 30.1300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.9300 0.0000 30.1300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.9300 0.0000 30.1300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[2]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 9.7240 54.6060 9.9240 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 9.7240 54.6060 9.9240 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 9.7240 54.6060 9.9240 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 9.7240 54.6060 9.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 9.7240 54.6060 9.9240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB1

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.7380 0.0000 24.9380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.7380 0.0000 24.9380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.7380 0.0000 24.9380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.7380 0.0000 24.9380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.7380 0.0000 24.9380 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.268128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.268128 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.2980 0.0000 31.4980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.2980 0.0000 31.4980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.2980 0.0000 31.4980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.2980 0.0000 31.4980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.2980 0.0000 31.4980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.6660 0.0000 32.8660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.6660 0.0000 32.8660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.6660 0.0000 32.8660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.6660 0.0000 32.8660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.6660 0.0000 32.8660 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I1[1]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.6010 0.0000 30.8010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.6010 0.0000 30.8010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.6010 0.0000 30.8010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.6010 0.0000 30.8010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.6010 0.0000 30.8010 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.268128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.268128 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8320 0.0000 34.0320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8320 0.0000 34.0320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8320 0.0000 34.0320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8320 0.0000 34.0320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8320 0.0000 34.0320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB1

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.6880 0.0000 22.8880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[3]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.3370 0.0000 33.5370 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.268308 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.268308 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.0950 0.0000 26.2950 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.267768 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.267768 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 132.5570 54.6060 132.7570 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 132.5570 54.6060 132.7570 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 132.5570 54.6060 132.7570 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 132.5570 54.6060 132.7570 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 132.5570 54.6060 132.7570 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 128.5670 54.6060 128.7670 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 128.5670 54.6060 128.7670 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 128.5670 54.6060 128.7670 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 128.5670 54.6060 128.7670 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 128.5670 54.6060 128.7670 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 132.5230 0.2000 132.7230 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 132.5230 0.2000 132.7230 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 132.5230 0.2000 132.7230 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 132.5230 0.2000 132.7230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS2

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 101.2310 54.6060 101.4310 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 101.2310 54.6060 101.4310 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 101.2310 54.6060 101.4310 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 101.2310 54.6060 101.4310 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 101.2310 54.6060 101.4310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[5]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 117.7010 54.6060 117.9010 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 117.7010 54.6060 117.9010 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 117.7010 54.6060 117.9010 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 117.7010 54.6060 117.9010 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 117.7010 54.6060 117.9010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[2]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 108.8790 54.6060 109.0790 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 108.8790 54.6060 109.0790 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 108.8790 54.6060 109.0790 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 108.8790 54.6060 109.0790 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 108.8790 54.6060 109.0790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[4]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 126.5180 54.6060 126.7180 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 126.5180 54.6060 126.7180 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 126.5180 54.6060 126.7180 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 126.5180 54.6060 126.7180 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 126.5180 54.6060 126.7180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 119.2880 54.6060 119.4880 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 119.2880 54.6060 119.4880 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 119.2880 54.6060 119.4880 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 119.2880 54.6060 119.4880 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 119.2880 54.6060 119.4880 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[1]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 25.9300 54.6060 26.1300 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 25.9300 54.6060 26.1300 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 25.9300 54.6060 26.1300 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 25.9300 54.6060 26.1300 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 25.9300 54.6060 26.1300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A1[6]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 126.5180 0.2000 126.7180 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 126.5180 0.2000 126.7180 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 126.5180 0.2000 126.7180 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 126.5180 0.2000 126.7180 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 126.5180 0.2000 126.7180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 119.2880 0.2000 119.4880 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 119.2880 0.2000 119.4880 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 119.2880 0.2000 119.4880 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 119.2880 0.2000 119.4880 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 119.2880 0.2000 119.4880 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 117.7010 0.2000 117.9010 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 117.7010 0.2000 117.9010 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 117.7010 0.2000 117.9010 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 117.7010 0.2000 117.9010 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 117.7010 0.2000 117.9010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 110.4680 0.2000 110.6680 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 110.4680 0.2000 110.6680 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 110.4680 0.2000 110.6680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 110.4680 0.2000 110.6680 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 110.4680 0.2000 110.6680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 108.8790 0.2000 109.0790 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 108.8790 0.2000 109.0790 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 108.8790 0.2000 109.0790 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 108.8790 0.2000 109.0790 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 108.8790 0.2000 109.0790 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[4]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 101.2310 0.2000 101.4310 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 101.2310 0.2000 101.4310 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 101.2310 0.2000 101.4310 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 101.2310 0.2000 101.4310 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 101.2310 0.2000 101.4310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.9300 0.2000 26.1300 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 25.9300 0.2000 26.1300 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 25.9300 0.2000 26.1300 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 25.9300 0.2000 26.1300 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 25.9300 0.2000 26.1300 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A2[6]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.7240 0.2000 9.9240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB2

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.2290 0.0000 29.4290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.2290 0.0000 29.4290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.2290 0.0000 29.4290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.2290 0.0000 29.4290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.2290 0.0000 29.4290 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.268308 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.268308 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.9650 0.0000 32.1650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.9650 0.0000 32.1650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.9650 0.0000 32.1650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.9650 0.0000 32.1650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.9650 0.0000 32.1650 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.268308 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.268308 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.0560 0.0000 24.2560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I2[2]

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 129.4130 54.6060 129.6130 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 129.4130 54.6060 129.6130 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 129.4130 54.6060 129.6130 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 129.4130 54.6060 129.6130 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 129.4130 54.6060 129.6130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.1170 0.2000 17.3170 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.4060 17.1570 54.6060 17.3570 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.1170 0.2000 17.3170 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 17.1570 54.6060 17.3570 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.1170 0.2000 17.3170 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 17.1570 54.6060 17.3570 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.1170 0.2000 17.3170 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 17.1570 54.6060 17.3570 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 17.1570 54.6060 17.3570 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE1

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.5280 139.4840 3.8280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.4290 139.4840 4.7280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.3280 139.4840 14.6280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.2290 139.4840 15.5290 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.4280 139.4840 49.7280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.3290 139.4840 50.6290 139.7840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.3590 0.0000 23.5590 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.267528 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.267528 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 0.8280 139.4840 1.1280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.7290 139.4840 2.0280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.6280 139.4840 11.9290 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.5290 139.4840 12.8280 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.0280 139.4840 53.3270 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.1290 139.4840 52.4290 139.7840 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 52.5790 139.4840 52.8790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.4780 139.4840 44.7770 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.6780 139.4840 42.9780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.5790 139.4840 43.8790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.1780 139.4840 47.4780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.6780 139.4840 51.9780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.4780 139.4840 53.7780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.2780 139.4840 46.5780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.0790 139.4840 48.3790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.9780 139.4840 49.2770 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.3790 139.4840 45.6800 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.8790 139.4840 50.1800 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.2780 139.4840 37.5780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.7780 139.4840 42.0780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.9780 139.4840 40.2770 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.1780 139.4840 38.4780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.0790 139.4840 39.3790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.5790 139.4840 34.8780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.8790 139.4840 41.1800 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.3780 139.4840 36.6790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.4780 139.4840 35.7790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.6790 139.4840 33.9780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.7790 139.4840 33.0790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.0790 139.4840 30.3780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.1790 139.4840 29.4780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.2790 139.4840 28.5790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.3780 139.4840 27.6780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.9780 139.4840 31.2790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.8780 139.4840 32.1790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.4790 139.4840 26.7790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.5780 139.4840 25.8780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.7790 139.4840 24.0780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.8790 139.4840 23.1790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.1790 139.4840 20.4790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.0780 139.4840 21.3780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.9780 139.4840 22.2790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.6780 139.4840 24.9790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.6780 139.4840 15.9780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.7790 139.4840 15.0780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.9790 139.4840 13.2790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.8780 139.4840 14.1780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.2790 139.4840 19.5790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.3780 139.4840 18.6790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.4780 139.4840 17.7790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.5780 139.4840 16.8790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.0780 139.4840 12.3780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.6790 139.4840 6.9780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.1790 139.4840 11.4780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.7790 139.4840 6.0790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.5790 139.4840 7.8780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.2790 139.4840 10.5790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.3780 139.4840 9.6790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.4780 139.4840 8.7790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.0780 139.4840 3.3780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.1790 139.4840 2.4790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.2780 139.4840 1.5780 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.8780 139.4840 5.1790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.9780 139.4840 4.2790 139.7840 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.7780 139.4840 51.0780 139.7840 ;
    END
  END VSS

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.4060 16.7390 54.6060 16.9390 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 16.7390 0.2000 16.9390 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.7390 0.2000 16.9390 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.4060 16.7390 54.6060 16.9390 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7390 0.2000 16.9390 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.4060 16.7390 54.6060 16.9390 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.7390 0.2000 16.9390 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.4060 16.7390 54.6060 16.9390 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.4060 16.7390 54.6060 16.9390 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB1
  OBS
    LAYER M3 ;
      RECT 0.0000 133.4570 54.6060 139.7840 ;
      RECT 0.0000 127.4180 53.7060 139.7840 ;
      RECT 0.0000 127.4180 53.7060 139.7840 ;
      RECT 0.0000 127.4180 53.7060 139.7840 ;
      RECT 0.0000 127.4180 53.7060 139.7840 ;
      RECT 0.0000 131.8570 53.7060 133.4570 ;
      RECT 0.0000 130.3130 53.7060 131.8570 ;
      RECT 0.0000 127.8670 53.7060 130.3130 ;
      RECT 0.0000 127.4180 53.7060 127.8670 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 125.8180 53.7060 127.4180 ;
      RECT 21.3000 0.0000 21.9880 0.9000 ;
      RECT 53.1050 130.3130 54.6060 131.8570 ;
      RECT 53.7060 127.4180 54.6060 127.8670 ;
      RECT 0.0000 120.1880 54.6060 125.8180 ;
      RECT 0.0000 111.3680 54.6060 117.0010 ;
      RECT 0.0000 102.1310 54.6060 108.1790 ;
      RECT 0.0000 26.8300 54.6060 100.5310 ;
      RECT 0.0000 18.0570 54.6060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 18.0570 ;
      RECT 0.0000 10.6240 54.6060 16.0390 ;
      RECT 0.0000 0.0000 19.7000 9.0240 ;
      RECT 0.0000 0.9000 54.6060 9.0240 ;
      RECT 0.0000 0.0000 19.7000 0.9000 ;
      RECT 0.9000 117.0010 53.7060 120.1880 ;
      RECT 0.9000 108.1790 53.7060 111.3680 ;
      RECT 0.9000 100.5310 53.7060 102.1310 ;
      RECT 0.9000 25.2300 53.7060 26.8300 ;
      RECT 0.9000 16.0390 53.7060 18.0170 ;
      RECT 0.9000 9.0240 53.7060 10.6240 ;
      RECT 34.7320 0.0000 54.6060 9.0240 ;
      RECT 34.7320 0.0000 54.6060 0.9000 ;
    LAYER M2 ;
      RECT 0.0000 127.4180 0.9000 128.6710 ;
      RECT 53.7060 127.4180 54.6060 127.8670 ;
      RECT 21.3000 0.0000 21.9880 0.9000 ;
      RECT 0.0000 130.2710 1.5010 131.8230 ;
      RECT 53.1050 130.3130 54.6060 131.8570 ;
      RECT 0.0000 120.1880 54.6060 125.8180 ;
      RECT 0.0000 111.3680 54.6060 117.0010 ;
      RECT 0.0000 102.1310 54.6060 108.1790 ;
      RECT 0.0000 26.8300 54.6060 100.5310 ;
      RECT 0.0000 18.0570 54.6060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 18.0570 ;
      RECT 0.0000 10.6240 54.6060 16.0390 ;
      RECT 0.0000 0.0000 19.7000 9.0240 ;
      RECT 0.0000 0.9000 54.6060 9.0240 ;
      RECT 0.0000 0.0000 19.7000 0.9000 ;
      RECT 0.9000 131.8230 53.7060 131.8570 ;
      RECT 0.9000 130.3130 53.7060 131.8230 ;
      RECT 0.9000 130.2710 53.7060 130.3130 ;
      RECT 0.9000 128.6710 53.7060 130.2710 ;
      RECT 0.9000 127.8670 53.7060 128.6710 ;
      RECT 0.9000 127.4180 53.7060 127.8670 ;
      RECT 0.9000 125.8180 53.7060 127.4180 ;
      RECT 0.9000 117.0010 53.7060 120.1880 ;
      RECT 0.9000 108.1790 53.7060 111.3680 ;
      RECT 0.9000 100.5310 53.7060 102.1310 ;
      RECT 0.9000 25.2300 53.7060 26.8300 ;
      RECT 0.9000 16.0390 53.7060 18.0170 ;
      RECT 0.9000 9.0240 53.7060 10.6240 ;
      RECT 34.7320 0.0000 54.6060 9.0240 ;
      RECT 34.7320 0.0000 54.6060 0.9000 ;
      RECT 0.0000 133.4570 54.6060 139.7840 ;
      RECT 0.0000 133.4230 53.7060 139.7840 ;
      RECT 0.0000 133.4230 53.7060 133.4570 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 131.8570 53.7060 133.4230 ;
    LAYER M1 ;
      RECT 0.0000 118.5010 0.8000 118.6880 ;
      RECT 53.8060 118.5010 54.6060 118.6880 ;
      RECT 0.0000 109.6790 54.6060 109.8680 ;
      RECT 53.8060 127.3180 54.6060 127.9670 ;
      RECT 21.2000 0.0000 22.0880 0.8000 ;
      RECT 0.0000 127.3180 0.8000 128.7710 ;
      RECT 0.0000 130.1710 1.5010 131.9230 ;
      RECT 0.0000 133.3230 53.8060 136.3240 ;
      RECT 53.1050 130.2130 54.6060 131.9570 ;
      RECT 0.8000 108.2790 53.8060 109.6790 ;
      RECT 0.8000 109.8680 53.8060 111.2800 ;
      RECT 0.8000 100.6310 53.8060 102.0310 ;
      RECT 0.0000 26.7300 54.6060 100.6310 ;
      RECT 0.0000 17.9570 54.6060 25.3300 ;
      RECT 0.0000 17.9170 53.8060 25.3300 ;
      RECT 0.0000 17.9170 53.8060 25.3300 ;
      RECT 0.0000 17.9170 53.8060 17.9570 ;
      RECT 0.8000 25.3300 53.8060 26.7300 ;
      RECT 0.8000 17.9570 53.8060 26.7300 ;
      RECT 0.8000 16.1390 53.8060 25.3300 ;
      RECT 0.8000 16.1390 53.8060 25.3300 ;
      RECT 0.8000 16.1390 53.8060 17.9170 ;
      RECT 0.0000 120.0880 54.6060 125.9180 ;
      RECT 0.0000 10.5240 54.6060 16.1390 ;
      RECT 0.0000 0.0000 19.8000 9.1240 ;
      RECT 0.0000 0.0000 19.8000 0.8000 ;
      RECT 0.0000 0.8000 54.6060 9.1240 ;
      RECT 0.8000 9.1240 53.8060 10.5240 ;
      RECT 0.8000 0.8000 53.8060 10.5240 ;
      RECT 34.6320 0.0000 54.6060 9.1240 ;
      RECT 34.6320 0.0000 54.6060 0.8000 ;
      RECT 0.8000 125.9180 53.8060 131.9230 ;
      RECT 0.8000 125.9180 53.8060 131.9230 ;
      RECT 0.8000 125.9180 53.8060 131.9230 ;
      RECT 0.8000 130.1710 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.8000 125.9180 53.8060 130.2130 ;
      RECT 0.0000 133.3570 54.6060 139.7840 ;
      RECT 0.8000 125.9180 53.8060 133.3230 ;
      RECT 0.8000 125.9180 53.8060 133.3230 ;
      RECT 0.8000 128.7710 53.8060 131.9570 ;
      RECT 0.8000 128.7710 53.8060 131.9570 ;
      RECT 0.8000 125.9180 53.8060 131.9570 ;
      RECT 0.0000 111.2680 54.6060 117.1010 ;
      RECT 0.0000 102.0310 54.6060 108.2790 ;
      RECT 0.8000 111.2680 53.8060 125.9180 ;
      RECT 0.8000 111.2680 53.8060 120.0880 ;
      RECT 0.8000 111.2680 53.8060 120.0880 ;
      RECT 0.8000 111.2680 53.8060 118.6880 ;
      RECT 0.8000 111.2680 53.8060 118.6880 ;
      RECT 0.8000 111.2680 53.8060 118.6880 ;
      RECT 0.8000 26.7300 53.8060 108.2790 ;
    LAYER PO ;
      RECT 0.0000 0.0000 54.6060 139.7840 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 54.6060 139.7840 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 54.6060 139.7840 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 54.6060 139.7840 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 54.6060 139.7840 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 54.6060 139.7840 ;
    LAYER M5 ;
      RECT 0.0000 138.7840 0.1280 139.7840 ;
      RECT 54.4780 138.7840 54.6060 139.7840 ;
      RECT 21.3000 0.0000 21.9880 0.9000 ;
      RECT 0.0000 130.2710 1.5010 131.8230 ;
      RECT 0.0000 127.4180 0.9000 128.6710 ;
      RECT 53.1050 130.3130 54.6060 131.8570 ;
      RECT 53.7060 127.4180 54.6060 127.8670 ;
      RECT 0.0000 120.1880 54.6060 125.8180 ;
      RECT 0.0000 111.3680 54.6060 117.0010 ;
      RECT 0.0000 102.1310 54.6060 108.1790 ;
      RECT 0.0000 26.8300 54.6060 100.5310 ;
      RECT 0.0000 18.0570 54.6060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 18.0570 ;
      RECT 0.0000 10.6240 54.6060 16.0390 ;
      RECT 0.0000 0.0000 19.7000 9.0240 ;
      RECT 0.0000 0.9000 54.6060 9.0240 ;
      RECT 0.0000 0.0000 19.7000 0.9000 ;
      RECT 0.9000 131.8230 53.7060 131.8570 ;
      RECT 0.9000 130.3130 53.7060 131.8230 ;
      RECT 0.9000 130.2710 53.7060 130.3130 ;
      RECT 0.9000 128.6710 53.7060 130.2710 ;
      RECT 0.9000 127.8670 53.7060 128.6710 ;
      RECT 0.9000 127.4180 53.7060 127.8670 ;
      RECT 0.9000 125.8180 53.7060 127.4180 ;
      RECT 0.9000 117.0010 53.7060 120.1880 ;
      RECT 0.9000 108.1790 53.7060 111.3680 ;
      RECT 0.9000 100.5310 53.7060 102.1310 ;
      RECT 0.9000 25.2300 53.7060 26.8300 ;
      RECT 0.9000 16.0390 53.7060 18.0170 ;
      RECT 0.9000 9.0240 53.7060 10.6240 ;
      RECT 34.7320 0.0000 54.6060 9.0240 ;
      RECT 34.7320 0.0000 54.6060 0.9000 ;
      RECT 0.0000 133.4570 54.6060 138.7840 ;
      RECT 0.0000 133.4230 53.7060 138.7840 ;
      RECT 0.0000 133.4230 53.7060 133.4570 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 0.9000 53.7060 138.7840 ;
      RECT 0.9000 131.8570 53.7060 133.4230 ;
    LAYER M4 ;
      RECT 21.3000 0.0000 21.9880 0.9000 ;
      RECT 0.0000 130.2710 1.5010 131.8230 ;
      RECT 0.0000 127.4180 0.9000 128.6710 ;
      RECT 53.1050 130.3130 54.6060 131.8570 ;
      RECT 53.7060 127.4180 54.6060 127.8670 ;
      RECT 0.0000 120.1880 54.6060 125.8180 ;
      RECT 0.0000 111.3680 54.6060 117.0010 ;
      RECT 0.0000 102.1310 54.6060 108.1790 ;
      RECT 0.0000 26.8300 54.6060 100.5310 ;
      RECT 0.0000 18.0570 54.6060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 25.2300 ;
      RECT 0.0000 18.0170 53.7060 18.0570 ;
      RECT 0.0000 10.6240 54.6060 16.0390 ;
      RECT 0.0000 0.0000 19.7000 9.0240 ;
      RECT 0.0000 0.9000 54.6060 9.0240 ;
      RECT 0.0000 0.0000 19.7000 0.9000 ;
      RECT 0.9000 131.8230 53.7060 131.8570 ;
      RECT 0.9000 130.3130 53.7060 131.8230 ;
      RECT 0.9000 130.2710 53.7060 130.3130 ;
      RECT 0.9000 128.6710 53.7060 130.2710 ;
      RECT 0.9000 127.8670 53.7060 128.6710 ;
      RECT 0.9000 127.4180 53.7060 127.8670 ;
      RECT 0.9000 125.8180 53.7060 127.4180 ;
      RECT 0.9000 117.0010 53.7060 120.1880 ;
      RECT 0.9000 108.1790 53.7060 111.3680 ;
      RECT 0.9000 100.5310 53.7060 102.1310 ;
      RECT 0.9000 25.2300 53.7060 26.8300 ;
      RECT 0.9000 16.0390 53.7060 18.0170 ;
      RECT 0.9000 9.0240 53.7060 10.6240 ;
      RECT 34.7320 0.0000 54.6060 9.0240 ;
      RECT 34.7320 0.0000 54.6060 0.9000 ;
      RECT 0.0000 133.4570 54.6060 139.7840 ;
      RECT 0.0000 133.4230 53.7060 139.7840 ;
      RECT 0.0000 133.4230 53.7060 133.4570 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 0.9000 53.7060 139.7840 ;
      RECT 0.9000 131.8570 53.7060 133.4230 ;
  END
END SRAMLP2RW128x4

MACRO SRAMLP2RW128x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 65.742 BY 141.691 ;
  SYMMETRY X Y R90 ;

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.2500 0.0000 36.4500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.2500 0.0000 36.4500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.2500 0.0000 36.4500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.2500 0.0000 36.4500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.2500 0.0000 36.4500 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279808 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279808 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.6170 0.0000 37.8170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.6170 0.0000 37.8170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.6170 0.0000 37.8170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.6170 0.0000 37.8170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.6170 0.0000 37.8170 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279748 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279748 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.9840 0.0000 39.1840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.9840 0.0000 39.1840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.9840 0.0000 39.1840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.9840 0.0000 39.1840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.9840 0.0000 39.1840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279808 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279808 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.3560 0.0000 40.5560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.3560 0.0000 40.5560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.3560 0.0000 40.5560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.3560 0.0000 40.5560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.3560 0.0000 40.5560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.280048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.280048 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.7240 0.0000 41.9240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.7240 0.0000 41.9240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.7240 0.0000 41.9240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.7240 0.0000 41.9240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.7240 0.0000 41.9240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.280048 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.280048 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.7900 0.0000 43.9900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.7900 0.0000 43.9900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.7900 0.0000 43.9900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.7900 0.0000 43.9900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.7900 0.0000 43.9900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.0930 0.0000 43.2930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.0930 0.0000 43.2930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.0930 0.0000 43.2930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.0930 0.0000 43.2930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.0930 0.0000 43.2930 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.280108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.280108 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.4610 0.0000 44.6610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.4610 0.0000 44.6610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.4610 0.0000 44.6610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.4610 0.0000 44.6610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.4610 0.0000 44.6610 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.280108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.280108 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.4220 0.0000 42.6220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.4220 0.0000 42.6220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.4220 0.0000 42.6220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.4220 0.0000 42.6220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.4220 0.0000 42.6220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.0540 0.0000 41.2540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.0540 0.0000 41.2540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.0540 0.0000 41.2540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.0540 0.0000 41.2540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.0540 0.0000 41.2540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.6860 0.0000 39.8860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.6860 0.0000 39.8860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.6860 0.0000 39.8860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.6860 0.0000 39.8860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.6860 0.0000 39.8860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.3180 0.0000 38.5180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.3180 0.0000 38.5180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.3180 0.0000 38.5180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.3180 0.0000 38.5180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.3180 0.0000 38.5180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.9500 0.0000 37.1500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.9500 0.0000 37.1500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.9500 0.0000 37.1500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.9500 0.0000 37.1500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.9500 0.0000 37.1500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.5820 0.0000 35.7820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.5820 0.0000 35.7820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.5820 0.0000 35.7820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.5820 0.0000 35.7820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.5820 0.0000 35.7820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.2140 0.0000 34.4140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.2140 0.0000 34.4140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.2140 0.0000 34.4140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.2140 0.0000 34.4140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.2140 0.0000 34.4140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4440 0.0000 32.6440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7080 0.0000 29.9080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3400 0.0000 28.5400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9720 0.0000 27.1720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 9.8930 65.7420 10.0930 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 9.8930 65.7420 10.0930 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 9.8930 65.7420 10.0930 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 9.8930 65.7420 10.0930 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 9.8930 65.7420 10.0930 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.16534 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16534 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.57204 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.57204 LAYER M2 ;
    ANTENNAMAXAREACAR 11.79836 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1582 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1582 LAYER M3 ;
    ANTENNAMAXAREACAR 12.88044 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1582 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1582 LAYER M4 ;
    ANTENNAMAXAREACAR 13.96244 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1582 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1582 LAYER M5 ;
    ANTENNAMAXAREACAR 15.04438 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4080 141.3900 60.7070 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.3080 141.3900 61.6070 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.0080 141.3900 19.3090 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.1090 141.3900 18.4090 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.5090 141.3900 5.8080 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.6090 141.3900 4.9080 141.6900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 253.2336 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 253.2336 LAYER M5 ;
  END VDDL

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.9550 0.0000 45.1550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.9550 0.0000 45.1550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.9550 0.0000 45.1550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.9550 0.0000 45.1550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.9550 0.0000 45.1550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.912217 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.912217 LAYER M2 ;
    ANTENNAMAXAREACAR 7.327361 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.38406 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.440691 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.49725 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB1

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5790 0.0000 20.7790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.903937 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.903937 LAYER M2 ;
    ANTENNAMAXAREACAR 7.26962 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.326324 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.382957 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.43952 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 134.9180 65.7420 135.1180 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 134.9180 65.7420 135.1180 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 134.9180 65.7420 135.1180 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 134.9180 65.7420 135.1180 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 134.9180 65.7420 135.1180 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.208245 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.208245 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.64293 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 30.68528 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.72744 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 131.4350 65.7420 131.6350 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 131.4350 65.7420 131.6350 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 131.4350 65.7420 131.6350 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 131.4350 65.7420 131.6350 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 131.4350 65.7420 131.6350 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
    ANTENNAGATEAREA 0.6282 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 4.021035 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.021035 LAYER M3 ;
    ANTENNAMAXAREACAR 14.30337 LAYER M3 ;
    ANTENNAGATEAREA 0.6282 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 14.54375 LAYER M4 ;
    ANTENNAGATEAREA 0.6282 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.78412 LAYER M5 ;
    ANTENNAGATEAREA 0.6282 LAYER M6 ;
    ANTENNAGATEAREA 0.6282 LAYER M7 ;
    ANTENNAGATEAREA 0.6282 LAYER M8 ;
    ANTENNAGATEAREA 0.6282 LAYER M9 ;
    ANTENNAGATEAREA 0.6282 LAYER MRDL ;
  END SD

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 131.7890 65.7420 131.9890 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 131.7890 65.7420 131.9890 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 131.7890 65.7420 131.9890 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 131.7890 65.7420 131.9890 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 131.7890 65.7420 131.9890 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END DS1

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 134.9340 0.2000 135.1340 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 134.9340 0.2000 135.1340 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 134.9340 0.2000 135.1340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 134.9340 0.2000 135.1340 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 134.9340 0.2000 135.1340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.208245 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.208245 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.010992 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.010992 LAYER M2 ;
    ANTENNAMAXAREACAR 22.26466 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1936 LAYER M3 ;
    ANTENNAMAXAREACAR 29.87695 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 2.4097 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4097 LAYER M4 ;
    ANTENNAMAXAREACAR 78.26437 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8940 0.2000 10.0940 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8940 0.2000 10.0940 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8940 0.2000 10.0940 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8940 0.2000 10.0940 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8940 0.2000 10.0940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15652 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15652 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56658 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56658 LAYER M2 ;
    ANTENNAMAXAREACAR 11.76099 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAMAXAREACAR 12.78964 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 13.81822 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 14.84674 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8680 0.0000 23.0680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2360 0.0000 24.4360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5220 0.0000 23.7220 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278968 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8990 0.0000 25.0990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8990 0.0000 25.0990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8990 0.0000 25.0990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8990 0.0000 25.0990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8990 0.0000 25.0990 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279028 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279028 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2690 0.0000 26.4690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2690 0.0000 26.4690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2690 0.0000 26.4690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2690 0.0000 26.4690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2690 0.0000 26.4690 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279628 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6380 0.0000 27.8380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6380 0.0000 27.8380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6380 0.0000 27.8380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6380 0.0000 27.8380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6380 0.0000 27.8380 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279688 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279688 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9920 0.0000 29.1920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9920 0.0000 29.1920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9920 0.0000 29.1920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9920 0.0000 29.1920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9920 0.0000 29.1920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.278848 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.278848 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7440 0.0000 31.9440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7440 0.0000 31.9440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7440 0.0000 31.9440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7440 0.0000 31.9440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7440 0.0000 31.9440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279928 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279928 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.5160 0.0000 33.7160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.5160 0.0000 33.7160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.5160 0.0000 33.7160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.5160 0.0000 33.7160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.5160 0.0000 33.7160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.304168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.304168 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.8850 0.0000 35.0850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.8850 0.0000 35.0850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.8850 0.0000 35.0850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.8850 0.0000 35.0850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.8850 0.0000 35.0850 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279988 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279988 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 103.8840 65.7420 104.0840 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 103.8840 65.7420 104.0840 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 103.8840 65.7420 104.0840 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 103.8840 65.7420 104.0840 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 103.8840 65.7420 104.0840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.285564 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.285564 LAYER M1 ;
    ANTENNAGATEAREA 20.0784 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 55.16673 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.16673 LAYER M2 ;
    ANTENNAMAXAREACAR 15.87503 LAYER M2 ;
    ANTENNAGATEAREA 20.4492 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 9.74912 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.74912 LAYER M3 ;
    ANTENNAMAXAREACAR 6.196228 LAYER M3 ;
    ANTENNAGATEAREA 20.4492 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 20.7688 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.7688 LAYER M4 ;
    ANTENNAMAXAREACAR 17.36739 LAYER M4 ;
    ANTENNAGATEAREA 20.4492 LAYER M5 ;
    ANTENNAGATEAREA 20.4492 LAYER M6 ;
    ANTENNAGATEAREA 20.4492 LAYER M7 ;
    ANTENNAGATEAREA 20.4492 LAYER M8 ;
    ANTENNAGATEAREA 20.4492 LAYER M9 ;
    ANTENNAGATEAREA 20.4492 LAYER MRDL ;
  END A1[5]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 112.7050 65.7420 112.9050 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 112.7050 65.7420 112.9050 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 112.7050 65.7420 112.9050 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 112.7050 65.7420 112.9050 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 112.7050 65.7420 112.9050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.285564 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.285564 LAYER M1 ;
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 111.2990 65.7420 111.4990 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 111.2990 65.7420 111.4990 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 111.2990 65.7420 111.4990 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 111.2990 65.7420 111.4990 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 111.2990 65.7420 111.4990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.285564 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.285564 LAYER M1 ;
  END A1[4]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 121.5260 65.7420 121.7260 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 121.5260 65.7420 121.7260 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 121.5260 65.7420 121.7260 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 121.5260 65.7420 121.7260 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 121.5260 65.7420 121.7260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.285564 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.285564 LAYER M1 ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 120.1190 65.7420 120.3190 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 120.1190 65.7420 120.3190 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 120.1190 65.7420 120.3190 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 120.1190 65.7420 120.3190 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 120.1190 65.7420 120.3190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.285564 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.285564 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72094 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72094 LAYER M2 ;
    ANTENNAMAXAREACAR 21.14282 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAMAXAREACAR 25.25071 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 29.35832 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 33.46566 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[2]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 128.9380 65.7420 129.1380 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 128.9380 65.7420 129.1380 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 128.9380 65.7420 129.1380 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 128.9380 65.7420 129.1380 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 128.9380 65.7420 129.1380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.285564 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.285564 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72106 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72106 LAYER M2 ;
    ANTENNAMAXAREACAR 21.1461 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAMAXAREACAR 25.25398 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 29.36159 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 33.46893 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A1[0]

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 131.7440 0.2000 131.9440 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 131.7440 0.2000 131.9440 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 131.7440 0.2000 131.9440 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 131.7440 0.2000 131.9440 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 131.7440 0.2000 131.9440 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.0213 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.226368 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.226368 LAYER M2 ;
    ANTENNAMAXAREACAR 12.55466 LAYER M2 ;
    ANTENNAGATEAREA 0.0912 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 4.792016 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.792016 LAYER M3 ;
    ANTENNAMAXAREACAR 56.39783 LAYER M3 ;
    ANTENNAGATEAREA 0.0912 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.3032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3032 LAYER M4 ;
    ANTENNAMAXAREACAR 68.42108 LAYER M4 ;
    ANTENNAGATEAREA 0.0912 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.3032 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3032 LAYER M5 ;
    ANTENNAMAXAREACAR 71.74339 LAYER M5 ;
    ANTENNAGATEAREA 0.0912 LAYER M6 ;
    ANTENNAGATEAREA 0.0912 LAYER M7 ;
    ANTENNAGATEAREA 0.0912 LAYER M8 ;
    ANTENNAGATEAREA 0.0912 LAYER M9 ;
    ANTENNAGATEAREA 0.0912 LAYER MRDL ;
  END DS2

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.1510 0.2000 28.3510 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 28.1510 0.2000 28.3510 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 28.1510 0.2000 28.3510 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 28.1510 0.2000 28.3510 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 28.1510 0.2000 28.3510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
    ANTENNAGATEAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.84532 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.84532 LAYER M2 ;
    ANTENNAMAXAREACAR 48.77866 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAMAXAREACAR 55.93732 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 63.09551 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 70.25322 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[6]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 103.8850 0.2000 104.0850 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 103.8850 0.2000 104.0850 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 103.8850 0.2000 104.0850 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 103.8850 0.2000 104.0850 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 103.8850 0.2000 104.0850 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
    ANTENNAGATEAREA 19.7844 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 48.43278 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 48.43278 LAYER M2 ;
    ANTENNAMAXAREACAR 15.29231 LAYER M2 ;
    ANTENNAGATEAREA 20.1552 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 11.04086 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.04086 LAYER M3 ;
    ANTENNAMAXAREACAR 6.267273 LAYER M3 ;
    ANTENNAGATEAREA 20.1552 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 8.7385 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7385 LAYER M4 ;
    ANTENNAMAXAREACAR 16.27363 LAYER M4 ;
    ANTENNAGATEAREA 49.2756 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 5408.045 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5408.045 LAYER M5 ;
    ANTENNAMAXAREACAR 196.7247 LAYER M5 ;
    ANTENNAGATEAREA 49.2756 LAYER M6 ;
    ANTENNAGATEAREA 49.2756 LAYER M7 ;
    ANTENNAGATEAREA 49.2756 LAYER M8 ;
    ANTENNAGATEAREA 49.2756 LAYER M9 ;
    ANTENNAGATEAREA 49.2756 LAYER MRDL ;
  END A2[5]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 128.9380 0.2000 129.1380 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 128.9380 0.2000 129.1380 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 128.9380 0.2000 129.1380 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 128.9380 0.2000 129.1380 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 128.9380 0.2000 129.1380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72112 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72112 LAYER M2 ;
    ANTENNAMAXAREACAR 21.14774 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAMAXAREACAR 25.25562 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 29.36323 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 33.47057 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 121.5250 0.2000 121.7250 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 121.5250 0.2000 121.7250 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 121.5250 0.2000 121.7250 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 121.5250 0.2000 121.7250 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 121.5250 0.2000 121.7250 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72118 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72118 LAYER M2 ;
    ANTENNAMAXAREACAR 21.14938 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAMAXAREACAR 25.25726 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 29.36487 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 33.47221 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 120.1190 0.2000 120.3190 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 120.1190 0.2000 120.3190 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 120.1190 0.2000 120.3190 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 120.1190 0.2000 120.3190 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 120.1190 0.2000 120.3190 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 112.7050 0.2000 112.9050 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 112.7050 0.2000 112.9050 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 112.7050 0.2000 112.9050 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 112.7050 0.2000 112.9050 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 112.7050 0.2000 112.9050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 111.2990 0.2000 111.4990 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 111.2990 0.2000 111.4990 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 111.2990 0.2000 111.4990 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 111.2990 0.2000 111.4990 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 111.2990 0.2000 111.4990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.287616 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.287616 LAYER M1 ;
  END A2[4]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4410 0.2000 17.6410 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4410 0.2000 17.6410 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4410 0.2000 17.6410 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4410 0.2000 17.6410 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4410 0.2000 17.6410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15652 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15652 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15652 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15652 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAGATEAREA 0.0894 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.31546 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.31546 LAYER M4 ;
    ANTENNAMAXAREACAR 6.447766 LAYER M4 ;
    ANTENNAGATEAREA 0.0894 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 8.129664 LAYER M5 ;
    ANTENNAGATEAREA 0.0894 LAYER M6 ;
    ANTENNAGATEAREA 0.0894 LAYER M7 ;
    ANTENNAGATEAREA 0.0894 LAYER M8 ;
    ANTENNAGATEAREA 0.0894 LAYER M9 ;
    ANTENNAGATEAREA 0.0894 LAYER MRDL ;
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9070 0.2000 17.1070 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.9070 0.2000 17.1070 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.9070 0.2000 17.1070 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9070 0.2000 17.1070 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.9070 0.2000 17.1070 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15652 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15652 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15652 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15652 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER M4 ;
    ANTENNAMAXAREACAR 13.54174 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 17.65013 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0760 0.0000 31.2760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3740 0.0000 30.5740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3740 0.0000 30.5740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3740 0.0000 30.5740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3740 0.0000 30.5740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3740 0.0000 30.5740 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.279688 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.279688 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6040 0.0000 25.8040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5470 28.1510 65.7420 28.3510 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5470 28.1510 65.7420 28.3510 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5470 28.1510 65.7420 28.3510 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5470 28.1510 65.7420 28.3510 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5470 28.1510 65.7420 28.3510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1543 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1543 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.22084 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22084 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.90202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.90202 LAYER M3 ;
    ANTENNAMAXAREACAR 52.7624 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M4 ;
    ANTENNAMAXAREACAR 59.9208 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 67.07872 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[6]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 17.3630 65.7420 17.5630 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 17.3630 65.7420 17.5630 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 17.3630 65.7420 17.5630 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 17.3630 65.7420 17.5630 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 17.3630 65.7420 17.5630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15418 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15418 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15418 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15418 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.29884 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.29884 LAYER M4 ;
    ANTENNAMAXAREACAR 13.1664 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 17.56318 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.5420 16.9010 65.7420 17.1010 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.5420 16.9010 65.7420 17.1010 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.5420 16.9010 65.7420 17.1010 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.5420 16.9010 65.7420 17.1010 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.5420 16.9010 65.7420 17.1010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15418 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15418 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15418 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15418 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.423949 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.423949 LAYER M4 ;
    ANTENNAMAXAREACAR 14.03661 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 18.14497 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 64.0070 141.3900 64.3060 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.1080 141.3900 63.4080 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.9080 141.3900 11.2090 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8080 141.3900 12.1090 141.6900 ;
    END
    ANTENNADIFFAREA 10.95167 LAYER M5 ;
    ANTENNADIFFAREA 10.95167 LAYER M6 ;
    ANTENNADIFFAREA 10.95167 LAYER M7 ;
    ANTENNADIFFAREA 10.95167 LAYER M8 ;
    ANTENNADIFFAREA 10.95167 LAYER M9 ;
    ANTENNADIFFAREA 10.95167 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 253.2342 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 253.2342 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 5.0580 141.3900 5.3590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3590 141.3900 11.6580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6580 141.3900 8.9590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5580 141.3900 9.8590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4580 141.3900 1.7580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3590 141.3900 2.6590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2580 141.3900 3.5580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4590 141.3900 10.7590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7590 141.3900 8.0580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8590 141.3900 7.1580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9590 141.3900 6.2590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5580 141.3900 18.8590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6580 141.3900 17.9590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7580 141.3900 17.0590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8580 141.3900 16.1580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9590 141.3900 15.2580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0580 141.3900 14.3580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1590 141.3900 13.4590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2580 141.3900 12.5580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8580 141.3900 25.1590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1580 141.3900 22.4590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9590 141.3900 24.2580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0590 141.3900 23.3590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4590 141.3900 19.7590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5580 141.3900 36.8590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3580 141.3900 38.6580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3580 141.3900 47.6580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1580 141.3900 49.4570 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2590 141.3900 48.5590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7590 141.3900 35.0580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8580 141.3900 43.1580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4580 141.3900 46.7580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0590 141.3900 50.3600 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2590 141.3900 39.5590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7590 141.3900 44.0590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5590 141.3900 45.8600 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6580 141.3900 44.9570 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1580 141.3900 40.4570 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9580 141.3900 42.2580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0590 141.3900 41.3600 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2590 141.3900 30.5580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0580 141.3900 32.3590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5580 141.3900 63.8580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9590 141.3900 60.2590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3590 141.3900 56.6590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7590 141.3900 53.0590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9580 141.3900 51.2580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4570 141.3900 64.7570 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6570 141.3900 62.9570 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7580 141.3900 62.0580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8580 141.3900 61.1580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0580 141.3900 59.3580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1580 141.3900 58.4580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2580 141.3900 57.5580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4580 141.3900 55.7580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5580 141.3900 54.8580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6580 141.3900 53.9580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8580 141.3900 52.1580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8590 141.3900 34.1580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9590 141.3900 33.2590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7580 141.3900 26.0580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1580 141.3900 31.4590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6590 141.3900 26.9590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4580 141.3900 37.7580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6580 141.3900 35.9590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5580 141.3900 27.8580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4590 141.3900 28.7590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3590 141.3900 29.6580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2580 141.3900 21.5580 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3590 141.3900 20.6590 141.6900 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.1580 141.3900 4.4590 141.6900 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0000 0.8000 64.9420 9.2940 ;
      RECT 0.0000 0.8000 64.9420 9.2940 ;
      RECT 0.0000 0.8000 65.7420 9.2930 ;
      RECT 45.7550 0.0000 65.7420 9.2930 ;
      RECT 45.7550 0.0000 65.7420 0.8000 ;
      RECT 0.8000 131.1440 64.9420 134.3180 ;
      RECT 0.8000 131.1440 64.9420 134.3180 ;
      RECT 0.8000 131.1440 64.9420 134.3180 ;
      RECT 0.8000 128.3380 64.9420 134.3180 ;
      RECT 0.8000 128.3380 64.9420 134.3180 ;
      RECT 0.8000 128.3380 64.9420 132.5890 ;
      RECT 0.8000 128.3380 64.9420 132.5890 ;
      RECT 0.8000 130.8350 64.9420 131.1440 ;
      RECT 0.0000 135.7340 65.7420 141.6910 ;
      RECT 0.8000 132.5890 64.9420 135.7340 ;
      RECT 0.8000 131.1440 64.9420 135.7340 ;
      RECT 0.8000 131.1440 64.9420 135.7340 ;
      RECT 0.8000 128.3380 64.9420 135.7340 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 131.1440 64.9420 135.7180 ;
      RECT 0.8000 128.3380 64.9420 135.7180 ;
      RECT 0.8000 128.3380 64.9420 135.7180 ;
      RECT 0.8000 128.3380 64.9420 135.7180 ;
      RECT 0.8000 128.3380 64.9420 135.7180 ;
      RECT 0.8000 128.3380 64.9420 135.7180 ;
      RECT 64.9420 129.7380 65.7420 130.8350 ;
      RECT 21.3790 0.0000 22.2680 0.8000 ;
      RECT 64.2410 132.5890 65.7420 134.3180 ;
      RECT 0.0000 129.7380 0.8000 131.1440 ;
      RECT 62.7410 135.7180 65.7420 135.7340 ;
      RECT 0.0000 132.5440 1.5010 134.3340 ;
      RECT 0.0000 0.0000 19.9790 9.2930 ;
      RECT 0.0000 0.0000 19.9790 0.8000 ;
      RECT 0.0000 122.3260 65.7420 128.3380 ;
      RECT 0.8000 9.2940 64.9420 10.6930 ;
      RECT 0.0000 18.2410 65.7420 27.5510 ;
      RECT 0.0000 16.3010 64.9420 16.3070 ;
      RECT 0.0000 10.6940 64.9420 16.3070 ;
      RECT 0.0000 10.6940 64.9420 16.3070 ;
      RECT 0.0000 10.6940 64.9420 16.3070 ;
      RECT 0.0000 10.6940 65.7420 16.3010 ;
      RECT 0.8000 18.1630 65.7420 27.5510 ;
      RECT 0.8000 18.1630 65.7420 27.5510 ;
      RECT 0.8000 18.1630 65.7420 27.5510 ;
      RECT 0.8000 10.6940 64.9420 27.5510 ;
      RECT 0.8000 10.6940 64.9420 27.5510 ;
      RECT 0.8000 10.6940 64.9420 27.5510 ;
      RECT 0.8000 18.1630 65.7420 18.2410 ;
      RECT 0.8000 16.3070 64.9420 18.1630 ;
      RECT 0.8000 10.6930 65.7420 16.3010 ;
      RECT 0.8000 10.6930 65.7420 16.3010 ;
      RECT 0.8000 10.6930 65.7420 16.3010 ;
      RECT 0.8000 9.2940 64.9420 16.3010 ;
      RECT 0.8000 9.2940 64.9420 16.3010 ;
      RECT 0.8000 9.2940 64.9420 16.3010 ;
      RECT 0.8000 10.6930 65.7420 10.6940 ;
      RECT 0.0000 122.3250 64.9420 122.3260 ;
      RECT 0.8000 119.5190 64.9420 122.3250 ;
      RECT 0.0000 113.5050 65.7420 119.5190 ;
      RECT 0.0000 104.6850 65.7420 110.6990 ;
      RECT 0.8000 113.5050 64.9420 122.3250 ;
      RECT 0.8000 113.5050 64.9420 122.3250 ;
      RECT 0.8000 110.6990 64.9420 113.5050 ;
      RECT 0.8000 104.6850 64.9420 113.5050 ;
      RECT 0.0000 103.2840 64.9420 103.2850 ;
      RECT 0.0000 28.9510 64.9420 103.2850 ;
      RECT 0.0000 28.9510 64.9420 103.2850 ;
      RECT 0.0000 28.9510 64.9420 103.2850 ;
      RECT 0.0000 28.9510 65.7420 103.2840 ;
      RECT 0.8000 104.6840 65.7420 104.6850 ;
      RECT 0.8000 103.2850 64.9420 104.6840 ;
      RECT 0.8000 28.9510 64.9420 104.6840 ;
      RECT 0.8000 28.9510 64.9420 104.6840 ;
      RECT 0.8000 28.9510 64.9420 104.6840 ;
      RECT 0.8000 27.5510 64.9470 103.2840 ;
      RECT 0.8000 27.5510 64.9470 28.9510 ;
      RECT 0.0000 9.2930 64.9420 9.2940 ;
      RECT 0.0000 0.8000 64.9420 9.2940 ;
    LAYER PO ;
      RECT 0.0000 0.0000 65.7420 141.6910 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 19.8790 9.1930 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 122.4260 65.7420 128.2380 ;
      RECT 0.9000 9.1940 64.8420 10.7930 ;
      RECT 0.0000 18.3410 65.7420 27.4510 ;
      RECT 0.0000 16.2010 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 65.7420 16.2010 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 18.3410 ;
      RECT 0.9000 16.2070 64.8420 18.2630 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 10.7940 ;
      RECT 0.0000 122.4250 64.8420 122.4260 ;
      RECT 0.0000 113.6050 65.7420 119.4190 ;
      RECT 0.9000 119.4190 64.8420 122.4250 ;
      RECT 0.9000 113.6050 64.8420 122.4250 ;
      RECT 0.0000 104.7850 65.7420 110.5990 ;
      RECT 0.9000 110.5990 64.8420 113.6050 ;
      RECT 0.0000 103.1840 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 65.7420 103.1840 ;
      RECT 0.9000 104.7840 65.7420 110.5990 ;
      RECT 0.9000 104.7840 65.7420 104.7850 ;
      RECT 0.9000 103.1850 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 27.4510 64.8470 103.1840 ;
      RECT 0.9000 27.4510 64.8470 29.0510 ;
      RECT 0.0000 9.1930 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 0.9000 ;
      RECT 0.9000 130.7350 64.8420 131.0440 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 132.6890 ;
      RECT 0.9000 128.2380 64.8420 132.6890 ;
      RECT 0.0000 135.8340 65.7420 141.6910 ;
      RECT 0.9000 132.6890 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8340 ;
      RECT 0.9000 128.2380 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 64.8420 129.8380 65.7420 130.7350 ;
      RECT 21.4790 0.0000 22.1680 0.9000 ;
      RECT 64.2410 132.6890 65.7420 134.2180 ;
      RECT 0.0000 132.6440 0.9000 132.6890 ;
      RECT 0.0000 129.8380 0.9000 131.0440 ;
      RECT 0.0000 132.6890 1.5010 134.2340 ;
      RECT 62.7410 135.8180 65.7420 135.8340 ;
    LAYER M4 ;
      RECT 0.0000 29.0510 65.7420 103.1840 ;
      RECT 0.9000 104.7840 65.7420 110.5990 ;
      RECT 0.9000 104.7840 65.7420 104.7850 ;
      RECT 0.9000 103.1850 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 27.4510 64.8470 103.1840 ;
      RECT 0.9000 27.4510 64.8470 29.0510 ;
      RECT 0.0000 9.1930 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 0.9000 ;
      RECT 0.9000 130.7350 64.8420 131.0440 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 132.6890 ;
      RECT 0.9000 128.2380 64.8420 132.6890 ;
      RECT 0.0000 135.8340 65.7420 141.6910 ;
      RECT 0.9000 132.6890 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8340 ;
      RECT 0.9000 128.2380 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 21.4790 0.0000 22.1680 0.9000 ;
      RECT 0.0000 132.6890 1.5010 134.2340 ;
      RECT 0.0000 129.8380 0.9000 131.0440 ;
      RECT 0.0000 132.6440 0.9000 132.6890 ;
      RECT 62.7410 135.8180 65.7420 135.8340 ;
      RECT 64.2410 132.6890 65.7420 134.2180 ;
      RECT 64.8420 129.8380 65.7420 130.7350 ;
      RECT 0.0000 0.0000 19.8790 9.1930 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 122.4260 65.7420 128.2380 ;
      RECT 0.9000 9.1940 64.8420 10.7930 ;
      RECT 0.0000 18.3410 65.7420 27.4510 ;
      RECT 0.0000 16.2010 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 65.7420 16.2010 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 18.3410 ;
      RECT 0.9000 16.2070 64.8420 18.2630 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 10.7940 ;
      RECT 0.0000 122.4250 64.8420 122.4260 ;
      RECT 0.0000 113.6050 65.7420 119.4190 ;
      RECT 0.9000 119.4190 64.8420 122.4250 ;
      RECT 0.9000 113.6050 64.8420 122.4250 ;
      RECT 0.0000 104.7850 65.7420 110.5990 ;
      RECT 0.9000 110.5990 64.8420 113.6050 ;
      RECT 0.0000 103.1840 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
    LAYER M3 ;
      RECT 21.4790 0.0000 22.1680 0.9000 ;
      RECT 0.0000 132.6890 1.5010 134.2340 ;
      RECT 0.0000 129.8380 0.9000 131.0440 ;
      RECT 0.0000 132.6440 0.9000 132.6890 ;
      RECT 62.7410 135.8180 65.7420 135.8340 ;
      RECT 64.2410 132.6890 65.7420 134.2180 ;
      RECT 64.8420 129.8380 65.7420 130.7350 ;
      RECT 0.0000 0.0000 19.8790 9.1930 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.0000 122.4260 65.7420 128.2380 ;
      RECT 0.9000 9.1940 64.8420 10.7930 ;
      RECT 0.0000 18.3410 65.7420 27.4510 ;
      RECT 0.0000 16.2010 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 65.7420 16.2010 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 18.3410 ;
      RECT 0.9000 16.2070 64.8420 18.2630 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 10.7940 ;
      RECT 0.0000 122.4250 64.8420 122.4260 ;
      RECT 0.0000 113.6050 65.7420 119.4190 ;
      RECT 0.9000 119.4190 64.8420 122.4250 ;
      RECT 0.9000 113.6050 64.8420 122.4250 ;
      RECT 0.0000 104.7850 65.7420 110.5990 ;
      RECT 0.9000 110.5990 64.8420 113.6050 ;
      RECT 0.0000 103.1840 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 65.7420 103.1840 ;
      RECT 0.9000 104.7840 65.7420 110.5990 ;
      RECT 0.9000 104.7840 65.7420 104.7850 ;
      RECT 0.9000 103.1850 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 27.4510 64.8470 103.1840 ;
      RECT 0.9000 27.4510 64.8470 29.0510 ;
      RECT 0.0000 9.1930 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 0.9000 ;
      RECT 0.9000 130.7350 64.8420 131.0440 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 132.6890 ;
      RECT 0.9000 128.2380 64.8420 132.6890 ;
      RECT 0.0000 135.8340 65.7420 141.6910 ;
      RECT 0.9000 132.6890 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8340 ;
      RECT 0.9000 128.2380 64.8420 135.8340 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 131.0440 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
      RECT 0.9000 128.2380 64.8420 135.8180 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 65.7420 141.6910 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 65.7420 141.6910 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 65.7420 141.6910 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 65.7420 141.6910 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 65.7420 141.6910 ;
    LAYER M5 ;
      RECT 65.4570 140.6900 65.7420 141.6910 ;
      RECT 0.0000 140.6900 0.7580 141.6910 ;
      RECT 21.4790 0.0000 22.1680 0.9000 ;
      RECT 0.0000 129.8380 0.9000 131.0440 ;
      RECT 0.0000 132.6440 0.9000 132.6890 ;
      RECT 0.0000 132.6890 1.5010 134.2180 ;
      RECT 0.0000 134.2180 0.9000 134.2340 ;
      RECT 64.2410 132.6890 65.7420 134.2180 ;
      RECT 64.8420 129.8380 65.7420 130.7350 ;
      RECT 0.0000 0.0000 19.8790 9.1930 ;
      RECT 0.0000 0.0000 19.8790 0.9000 ;
      RECT 0.9000 130.7350 64.8420 131.0440 ;
      RECT 0.9000 18.2630 65.7420 18.3410 ;
      RECT 0.9000 16.2070 64.8420 18.2630 ;
      RECT 0.0000 18.3410 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.9000 18.2630 65.7420 27.4510 ;
      RECT 0.0000 16.2010 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 64.8420 16.2070 ;
      RECT 0.0000 10.7940 65.7420 16.2010 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7940 64.8420 27.4510 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 9.1940 64.8420 16.2010 ;
      RECT 0.9000 10.7930 65.7420 10.7940 ;
      RECT 0.9000 9.1940 64.8420 10.7930 ;
      RECT 0.0000 135.8340 65.7420 140.6900 ;
      RECT 0.9000 135.8180 65.7420 135.8340 ;
      RECT 0.9000 132.6890 64.8420 135.8340 ;
      RECT 0.9000 134.2180 64.8420 134.2340 ;
      RECT 0.9000 132.6890 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 131.0440 64.8420 134.2180 ;
      RECT 0.9000 130.7350 64.8420 134.2180 ;
      RECT 0.9000 129.8380 64.8420 134.2180 ;
      RECT 0.9000 130.7350 64.8420 134.2180 ;
      RECT 0.9000 129.8380 64.8420 134.2180 ;
      RECT 0.9000 130.7350 64.8420 134.2180 ;
      RECT 0.9000 129.8380 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 134.2180 ;
      RECT 0.9000 128.2380 64.8420 134.2180 ;
      RECT 0.0000 122.4260 65.7420 128.2380 ;
      RECT 0.0000 122.4250 64.8420 122.4260 ;
      RECT 0.0000 113.6050 65.7420 119.4190 ;
      RECT 0.9000 113.6050 64.8420 122.4260 ;
      RECT 0.9000 119.4190 64.8420 122.4250 ;
      RECT 0.0000 103.1840 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 64.8420 103.1850 ;
      RECT 0.0000 29.0510 65.7420 103.1840 ;
      RECT 0.9000 27.4510 64.8470 103.1840 ;
      RECT 0.9000 27.4510 64.8470 29.0510 ;
      RECT 0.0000 104.7850 65.7420 110.5990 ;
      RECT 0.9000 110.5990 64.8420 113.6050 ;
      RECT 0.9000 104.7840 65.7420 110.5990 ;
      RECT 0.9000 104.7840 65.7420 104.7850 ;
      RECT 0.9000 103.1850 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.9000 29.0510 64.8420 104.7840 ;
      RECT 0.0000 9.1930 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 64.8420 9.1940 ;
      RECT 0.0000 0.9000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 9.1930 ;
      RECT 45.8550 0.0000 65.7420 0.9000 ;
  END
END SRAMLP2RW128x8

MACRO SRAMLP2RW128x16
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 87.63 BY 146.025 ;
  SYMMETRY X Y R90 ;

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 115.4320 87.6300 115.6320 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 115.4320 87.6300 115.6320 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 115.4320 87.6300 115.6320 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 115.4320 87.6300 115.6320 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 115.4320 87.6300 115.6320 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2887 LAYER M1 ;
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 108.2040 87.6300 108.4040 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 108.2040 87.6300 108.4040 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 108.2040 87.6300 108.4040 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 108.2040 87.6300 108.4040 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 108.2040 87.6300 108.4040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2887 LAYER M1 ;
    ANTENNAGATEAREA 1.098 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 6.23156 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.23156 LAYER M2 ;
    ANTENNAMAXAREACAR 13.72651 LAYER M2 ;
    ANTENNAGATEAREA 1.098 LAYER M3 ;
    ANTENNAGATEAREA 1.098 LAYER M4 ;
    ANTENNAGATEAREA 1.098 LAYER M5 ;
    ANTENNAGATEAREA 1.098 LAYER M6 ;
    ANTENNAGATEAREA 1.098 LAYER M7 ;
    ANTENNAGATEAREA 1.098 LAYER M8 ;
    ANTENNAGATEAREA 1.098 LAYER M9 ;
    ANTENNAGATEAREA 1.098 LAYER MRDL ;
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 32.4380 87.6300 32.6380 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 32.4380 87.6300 32.6380 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 32.4380 87.6300 32.6380 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 32.4380 87.6300 32.6380 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 32.4380 87.6300 32.6380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.23116 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23116 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.90322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.90322 LAYER M3 ;
    ANTENNAMAXAREACAR 52.67027 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 59.88584 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 67.10094 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[6]

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 139.2950 0.2000 139.4950 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 139.2950 0.2000 139.4950 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 139.2950 0.2000 139.4950 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 139.2950 0.2000 139.4950 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 139.2950 0.2000 139.4950 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.220395 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.220395 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.97487 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.0172 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.05933 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.3680 0.2000 17.5680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15256 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15256 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15256 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0894 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30916 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30916 LAYER M4 ;
    ANTENNAMAXAREACAR 6.377295 LAYER M4 ;
    ANTENNAGATEAREA 0.0894 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.072623 LAYER M5 ;
    ANTENNAGATEAREA 0.0894 LAYER M6 ;
    ANTENNAGATEAREA 0.0894 LAYER M7 ;
    ANTENNAGATEAREA 0.0894 LAYER M8 ;
    ANTENNAGATEAREA 0.0894 LAYER M9 ;
    ANTENNAGATEAREA 0.0894 LAYER MRDL ;
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.8340 0.2000 17.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15256 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15256 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15256 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.40684 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40684 LAYER M4 ;
    ANTENNAMAXAREACAR 13.56469 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.70587 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 133.1320 0.2000 133.3320 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 133.1320 0.2000 133.3320 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 133.1320 0.2000 133.3320 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 133.1320 0.2000 133.3320 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 133.1320 0.2000 133.3320 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288136 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288136 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.71716 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.71716 LAYER M2 ;
    ANTENNAMAXAREACAR 21.01074 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.15144 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.29185 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.432 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 125.8350 0.2000 126.0350 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 125.8350 0.2000 126.0350 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 125.8350 0.2000 126.0350 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 125.8350 0.2000 126.0350 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 125.8350 0.2000 126.0350 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288136 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288136 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.71716 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.71716 LAYER M2 ;
    ANTENNAMAXAREACAR 20.9955 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.13619 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.27661 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.41676 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 124.3140 0.2000 124.5140 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 124.3140 0.2000 124.5140 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 124.3140 0.2000 124.5140 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 124.3140 0.2000 124.5140 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 124.3140 0.2000 124.5140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288136 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288136 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.71716 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.71716 LAYER M2 ;
    ANTENNAMAXAREACAR 21.01413 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.15482 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.29524 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.43539 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 117.0000 0.2000 117.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 117.0000 0.2000 117.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 117.0000 0.2000 117.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 117.0000 0.2000 117.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 117.0000 0.2000 117.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288136 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288136 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.71716 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.71716 LAYER M2 ;
    ANTENNAMAXAREACAR 21.02091 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.1616 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.30202 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.44216 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 115.4820 0.2000 115.6820 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 115.4820 0.2000 115.6820 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 115.4820 0.2000 115.6820 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 115.4820 0.2000 115.6820 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 115.4820 0.2000 115.6820 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288136 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288136 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.71716 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.71716 LAYER M2 ;
    ANTENNAMAXAREACAR 20.9938 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.1345 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.27492 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.41506 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[4]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 133.0920 87.6300 133.2920 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 133.0920 87.6300 133.2920 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 133.0920 87.6300 133.2920 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 133.0920 87.6300 133.2920 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 133.0920 87.6300 133.2920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2887 LAYER M1 ;
  END A1[0]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 16.8280 87.6300 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 16.8280 87.6300 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 16.8280 87.6300 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 16.8280 87.6300 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 16.8280 87.6300 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.424789 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.424789 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END CSB1

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 17.2900 87.6300 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 17.2900 87.6300 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 17.2900 87.6300 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 17.2900 87.6300 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 17.2900 87.6300 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.29968 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.29968 LAYER M4 ;
    ANTENNAMAXAREACAR 13.19096 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.62284 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 1.0080 145.7250 1.3070 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9070 145.7250 2.2080 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.9100 145.7250 11.2090 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8090 145.7250 12.1100 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.7080 145.7250 85.0070 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.6070 145.7250 85.9080 146.0250 ;
    END
    ANTENNADIFFAREA 10.95167 LAYER M5 ;
    ANTENNADIFFAREA 10.95167 LAYER M6 ;
    ANTENNADIFFAREA 10.95167 LAYER M7 ;
    ANTENNADIFFAREA 10.95167 LAYER M8 ;
    ANTENNADIFFAREA 10.95167 LAYER M9 ;
    ANTENNADIFFAREA 10.95167 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 261.1671 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 261.1671 LAYER M5 ;
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 5.0580 145.7250 5.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9580 145.7250 60.2580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.1590 145.7250 4.4590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0570 145.7250 59.3570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2580 145.7250 3.5580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2580 145.7250 57.5570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4590 145.7250 1.7580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4580 145.7250 64.7570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6590 145.7250 8.9580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5580 145.7250 63.8580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7590 145.7250 8.0590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5590 145.7250 54.8590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7580 145.7250 53.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3580 145.7250 56.6580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4580 145.7250 55.7580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6580 145.7250 53.9580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3580 145.7250 65.6570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5590 145.7250 9.8580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1570 145.7250 67.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3580 145.7250 11.6590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2570 145.7250 66.5580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4580 145.7250 10.7590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3570 145.7250 74.6580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5580 145.7250 18.8590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0580 145.7250 68.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2590 145.7250 12.5590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8570 145.7250 70.1570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0580 145.7250 14.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9580 145.7250 69.2570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1590 145.7250 13.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4570 145.7250 73.7570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6580 145.7250 17.9580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5580 145.7250 72.8570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7590 145.7250 17.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7580 145.7250 71.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9590 145.7250 15.2590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6570 145.7250 71.9570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8580 145.7250 16.1580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2570 145.7250 75.5580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4580 145.7250 19.7590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1570 145.7250 76.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3580 145.7250 20.6590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7570 145.7250 80.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9580 145.7250 24.2590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4570 145.7250 82.7580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6580 145.7250 26.9590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.0580 145.7250 77.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2590 145.7250 21.5590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9580 145.7250 78.2580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1590 145.7250 22.4590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5580 145.7250 81.8570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7590 145.7250 26.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8570 145.7250 79.1570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0580 145.7250 23.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6580 145.7250 80.9580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8590 145.7250 25.1590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2580 145.7250 84.5580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4590 145.7250 28.7590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3570 145.7250 83.6570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5580 145.7250 27.8580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1570 145.7250 85.4570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3580 145.7250 29.6580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0580 145.7250 86.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2590 145.7250 30.5590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1590 145.7250 31.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9580 145.7250 33.2590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3580 145.7250 38.6590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4580 145.7250 37.7590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8580 145.7250 34.1590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0590 145.7250 32.3580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0590 145.7250 41.3590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5590 145.7250 36.8580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2580 145.7250 39.5580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6590 145.7250 35.9580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7590 145.7250 35.0590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9580 145.7250 42.2570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1580 145.7250 40.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8590 145.7250 43.1600 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8590 145.7250 52.1600 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3590 145.7250 47.6600 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7580 145.7250 44.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9580 145.7250 51.2570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6580 145.7250 44.9580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4580 145.7250 46.7570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2580 145.7250 48.5580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0590 145.7250 50.3590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1580 145.7250 49.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5590 145.7250 45.8590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8570 145.7250 61.1570 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3580 145.7250 2.6590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1570 145.7250 58.4580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9580 145.7250 6.2590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7570 145.7250 62.0580 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8580 145.7250 7.1590 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6570 145.7250 62.9580 146.0250 ;
    END
  END VSS

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.2070 0.0000 60.4070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.2070 0.0000 60.4070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.2070 0.0000 60.4070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.2070 0.0000 60.4070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.2070 0.0000 60.4070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.5240 0.0000 59.7240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.5240 0.0000 59.7240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.5240 0.0000 59.7240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.5240 0.0000 59.7240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.5240 0.0000 59.7240 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.8390 0.0000 59.0390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.8390 0.0000 59.0390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.8390 0.0000 59.0390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.8390 0.0000 59.0390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.8390 0.0000 59.0390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.1560 0.0000 58.3560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.1560 0.0000 58.3560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.1560 0.0000 58.3560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.1560 0.0000 58.3560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.1560 0.0000 58.3560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.3640 0.0000 66.5640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.3640 0.0000 66.5640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.3640 0.0000 66.5640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.3640 0.0000 66.5640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.3640 0.0000 66.5640 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[3]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.6790 0.0000 65.8790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.6790 0.0000 65.8790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.6790 0.0000 65.8790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.6790 0.0000 65.8790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.6790 0.0000 65.8790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.9960 0.0000 65.1960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.9960 0.0000 65.1960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.9960 0.0000 65.1960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.9960 0.0000 65.1960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.9960 0.0000 65.1960 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[10]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.3110 0.0000 64.5110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.3110 0.0000 64.5110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.3110 0.0000 64.5110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.3110 0.0000 64.5110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.3110 0.0000 64.5110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.6280 0.0000 63.8280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.6280 0.0000 63.8280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.6280 0.0000 63.8280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.6280 0.0000 63.8280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.6280 0.0000 63.8280 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.9430 0.0000 63.1430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.9430 0.0000 63.1430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.9430 0.0000 63.1430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.9430 0.0000 63.1430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.9430 0.0000 63.1430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 9.8200 87.6300 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 9.8200 87.6300 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 9.8200 87.6300 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 9.8200 87.6300 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 9.8200 87.6300 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15724 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15724 LAYER M1 ;
  END WEB1

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8210 0.2000 10.0210 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15256 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15256 LAYER M1 ;
    ANTENNAGATEAREA 18.7377 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 121.896 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 121.896 LAYER M2 ;
    ANTENNAMAXAREACAR 42.06476 LAYER M2 ;
    ANTENNAGATEAREA 29.3091 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 35.46363 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.46363 LAYER M3 ;
    ANTENNAMAXAREACAR 11.42129 LAYER M3 ;
    ANTENNAGATEAREA 29.3091 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 185.8102 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 185.8102 LAYER M4 ;
    ANTENNAMAXAREACAR 49.61441 LAYER M4 ;
    ANTENNAGATEAREA 29.3559 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 7536.405 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 7536.405 LAYER M5 ;
    ANTENNAMAXAREACAR 343.6991 LAYER M5 ;
    ANTENNAGATEAREA 29.3559 LAYER M6 ;
    ANTENNAGATEAREA 29.3559 LAYER M7 ;
    ANTENNAGATEAREA 29.3559 LAYER M8 ;
    ANTENNAGATEAREA 29.3559 LAYER M9 ;
    ANTENNAGATEAREA 29.3559 LAYER MRDL ;
  END WEB2

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 136.0520 0.2000 136.2520 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 136.0520 0.2000 136.2520 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 136.0520 0.2000 136.2520 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 136.0520 0.2000 136.2520 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 136.0520 0.2000 136.2520 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.2256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.381546 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.381546 LAYER M2 ;
    ANTENNAMAXAREACAR 6.268031 LAYER M2 ;
    ANTENNAGATEAREA 0.7194 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 11.08991 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.08991 LAYER M3 ;
    ANTENNAMAXAREACAR 23.318 LAYER M3 ;
    ANTENNAGATEAREA 0.7194 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4548 LAYER M4 ;
    ANTENNAMAXAREACAR 23.94968 LAYER M4 ;
    ANTENNAGATEAREA 0.7194 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4548 LAYER M5 ;
    ANTENNAMAXAREACAR 24.58135 LAYER M5 ;
    ANTENNAGATEAREA 0.7194 LAYER M6 ;
    ANTENNAGATEAREA 0.7194 LAYER M7 ;
    ANTENNAGATEAREA 0.7194 LAYER M8 ;
    ANTENNAGATEAREA 0.7194 LAYER M9 ;
    ANTENNAGATEAREA 0.7194 LAYER MRDL ;
  END DS2

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 136.0160 87.6300 136.2160 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 136.0160 87.6300 136.2160 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 136.0160 87.6300 136.2160 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 136.0160 87.6300 136.2160 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 136.0160 87.6300 136.2160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END DS1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 135.6620 87.6300 135.8620 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 135.6620 87.6300 135.8620 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 135.6620 87.6300 135.8620 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 135.6620 87.6300 135.8620 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 135.6620 87.6300 135.8620 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END SD

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.2100 145.7250 8.5090 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.1090 145.7250 9.4100 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.4090 145.7250 15.7080 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.3080 145.7250 16.6090 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.9080 145.7250 83.2070 146.0250 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.8070 145.7250 84.1080 146.0250 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 261.1671 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 261.1671 LAYER M5 ;
  END VDDL

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5800 0.0000 20.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5800 0.0000 20.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5800 0.0000 20.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5800 0.0000 20.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5800 0.0000 20.7800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.2682 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.55626 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.55626 LAYER M2 ;
    ANTENNAMAXAREACAR 6.76863 LAYER M2 ;
    ANTENNAGATEAREA 0.2682 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 7.333433 LAYER M3 ;
    ANTENNAGATEAREA 0.2682 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.898199 LAYER M4 ;
    ANTENNAGATEAREA 0.2682 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.462928 LAYER M5 ;
    ANTENNAGATEAREA 0.2682 LAYER M6 ;
    ANTENNAGATEAREA 0.2682 LAYER M7 ;
    ANTENNAGATEAREA 0.2682 LAYER M8 ;
    ANTENNAGATEAREA 0.2682 LAYER M9 ;
    ANTENNAGATEAREA 0.2682 LAYER MRDL ;
  END OEB2

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 139.2230 87.6300 139.4230 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 139.2230 87.6300 139.4230 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 139.2230 87.6300 139.4230 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 139.2230 87.6300 139.4230 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 139.2230 87.6300 139.4230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.238615 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.238615 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 28.47265 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.51495 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.55704 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.8440 0.0000 67.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.8440 0.0000 67.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.8440 0.0000 67.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.8440 0.0000 67.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.8440 0.0000 67.0440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.2682 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56214 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56214 LAYER M2 ;
    ANTENNAMAXAREACAR 6.790553 LAYER M2 ;
    ANTENNAGATEAREA 0.2682 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 7.355355 LAYER M3 ;
    ANTENNAGATEAREA 0.2682 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.92012 LAYER M4 ;
    ANTENNAGATEAREA 0.2682 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.484847 LAYER M5 ;
    ANTENNAGATEAREA 0.2682 LAYER M6 ;
    ANTENNAGATEAREA 0.2682 LAYER M7 ;
    ANTENNAGATEAREA 0.2682 LAYER M8 ;
    ANTENNAGATEAREA 0.2682 LAYER M9 ;
    ANTENNAGATEAREA 0.2682 LAYER MRDL ;
  END OEB1

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.8440 0.0000 46.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.8440 0.0000 46.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.8440 0.0000 46.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.8440 0.0000 46.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.8440 0.0000 46.0440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.1590 0.0000 45.3590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.1590 0.0000 45.3590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.1590 0.0000 45.3590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.1590 0.0000 45.3590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.1590 0.0000 45.3590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0760 0.0000 44.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0760 0.0000 44.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0760 0.0000 44.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0760 0.0000 44.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0760 0.0000 44.2760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.3670 0.0000 53.5670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.3670 0.0000 53.5670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.3670 0.0000 53.5670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.3670 0.0000 53.5670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.3670 0.0000 53.5670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.6840 0.0000 52.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.6840 0.0000 52.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.6840 0.0000 52.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.6840 0.0000 52.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.6840 0.0000 52.8840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.9990 0.0000 52.1990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.9990 0.0000 52.1990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.9990 0.0000 52.1990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.9990 0.0000 52.1990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.9990 0.0000 52.1990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.3160 0.0000 51.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.3160 0.0000 51.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.3160 0.0000 51.5160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.3160 0.0000 51.5160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.3160 0.0000 51.5160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.6310 0.0000 50.8310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.6310 0.0000 50.8310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.6310 0.0000 50.8310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.6310 0.0000 50.8310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.6310 0.0000 50.8310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.9480 0.0000 50.1480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.9480 0.0000 50.1480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.9480 0.0000 50.1480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.9480 0.0000 50.1480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.9480 0.0000 50.1480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.2630 0.0000 49.4630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.2630 0.0000 49.4630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.2630 0.0000 49.4630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.2630 0.0000 49.4630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.2630 0.0000 49.4630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.4710 0.0000 57.6710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.4710 0.0000 57.6710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.4710 0.0000 57.6710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.4710 0.0000 57.6710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.4710 0.0000 57.6710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.7880 0.0000 56.9880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.7880 0.0000 56.9880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.7880 0.0000 56.9880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.7880 0.0000 56.9880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.7880 0.0000 56.9880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.1030 0.0000 56.3030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.1030 0.0000 56.3030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.1030 0.0000 56.3030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.1030 0.0000 56.3030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.1030 0.0000 56.3030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.4200 0.0000 55.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.4200 0.0000 55.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.4200 0.0000 55.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.4200 0.0000 55.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.4200 0.0000 55.6200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.7350 0.0000 54.9350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.7350 0.0000 54.9350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.7350 0.0000 54.9350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.7350 0.0000 54.9350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.7350 0.0000 54.9350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.0520 0.0000 54.2520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.0520 0.0000 54.2520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.0520 0.0000 54.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.0520 0.0000 54.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.0520 0.0000 54.2520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.2600 0.0000 62.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.2600 0.0000 62.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.2600 0.0000 62.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.2600 0.0000 62.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.2600 0.0000 62.4600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[9]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.5750 0.0000 61.7750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.5750 0.0000 61.7750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.5750 0.0000 61.7750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.5750 0.0000 61.7750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.5750 0.0000 61.7750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.8920 0.0000 61.0920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.8920 0.0000 61.0920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.8920 0.0000 61.0920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.8920 0.0000 61.0920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.8920 0.0000 61.0920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O1[14]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.2340 0.0000 37.4340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.2340 0.0000 37.4340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.2340 0.0000 37.4340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.2340 0.0000 37.4340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.2340 0.0000 37.4340 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5490 0.0000 36.7490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5490 0.0000 36.7490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5490 0.0000 36.7490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5490 0.0000 36.7490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5490 0.0000 36.7490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8660 0.0000 36.0660 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8660 0.0000 36.0660 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8660 0.0000 36.0660 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8660 0.0000 36.0660 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8660 0.0000 36.0660 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1810 0.0000 35.3810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1810 0.0000 35.3810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1810 0.0000 35.3810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1810 0.0000 35.3810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1810 0.0000 35.3810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4980 0.0000 34.6980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4980 0.0000 34.6980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4980 0.0000 34.6980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4980 0.0000 34.6980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4980 0.0000 34.6980 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9170 0.0000 38.1170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9170 0.0000 38.1170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9170 0.0000 38.1170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9170 0.0000 38.1170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9170 0.0000 38.1170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9700 0.0000 40.1700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9700 0.0000 40.1700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9700 0.0000 40.1700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9700 0.0000 40.1700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9700 0.0000 40.1700 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2850 0.0000 39.4850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2850 0.0000 39.4850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2850 0.0000 39.4850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2850 0.0000 39.4850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2850 0.0000 39.4850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.6020 0.0000 38.8020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.6020 0.0000 38.8020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.6020 0.0000 38.8020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.6020 0.0000 38.8020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.6020 0.0000 38.8020 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3890 0.0000 43.5890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3890 0.0000 43.5890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3890 0.0000 43.5890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3890 0.0000 43.5890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3890 0.0000 43.5890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.7060 0.0000 42.9060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.7060 0.0000 42.9060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.7060 0.0000 42.9060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.7060 0.0000 42.9060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.7060 0.0000 42.9060 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0210 0.0000 42.2210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0210 0.0000 42.2210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0210 0.0000 42.2210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0210 0.0000 42.2210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0210 0.0000 42.2210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.3380 0.0000 41.5380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.3380 0.0000 41.5380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.3380 0.0000 41.5380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.3380 0.0000 41.5380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.3380 0.0000 41.5380 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6530 0.0000 40.8530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6530 0.0000 40.8530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6530 0.0000 40.8530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6530 0.0000 40.8530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6530 0.0000 40.8530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.5800 0.0000 48.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.5800 0.0000 48.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.5800 0.0000 48.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.5800 0.0000 48.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.5800 0.0000 48.7800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.8950 0.0000 48.0950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.8950 0.0000 48.0950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.8950 0.0000 48.0950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.8950 0.0000 48.0950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.8950 0.0000 48.0950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.2120 0.0000 47.4120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.2120 0.0000 47.4120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.2120 0.0000 47.4120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.2120 0.0000 47.4120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.2120 0.0000 47.4120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.5270 0.0000 46.7270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.5270 0.0000 46.7270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.5270 0.0000 46.7270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.5270 0.0000 46.7270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.5270 0.0000 46.7270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 108.1960 0.2000 108.3960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 108.1960 0.2000 108.3960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 108.1960 0.2000 108.3960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 108.1960 0.2000 108.3960 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 108.1960 0.2000 108.3960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288136 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288136 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.71716 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.71716 LAYER M2 ;
    ANTENNAMAXAREACAR 20.9938 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.1345 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.27492 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.41506 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.4400 0.2000 32.6400 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 32.4400 0.2000 32.6400 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 32.4400 0.2000 32.6400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.4400 0.2000 32.6400 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 32.4400 0.2000 32.6400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.273576 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.273576 LAYER M1 ;
    ANTENNAGATEAREA 0.309 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 8.4472 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.4472 LAYER M2 ;
    ANTENNAMAXAREACAR 38.32599 LAYER M2 ;
    ANTENNAGATEAREA 0.309 LAYER M3 ;
    ANTENNAGATEAREA 0.309 LAYER M4 ;
    ANTENNAGATEAREA 0.309 LAYER M5 ;
    ANTENNAGATEAREA 0.309 LAYER M6 ;
    ANTENNAGATEAREA 0.309 LAYER M7 ;
    ANTENNAGATEAREA 0.309 LAYER M8 ;
    ANTENNAGATEAREA 0.309 LAYER M9 ;
    ANTENNAGATEAREA 0.309 LAYER MRDL ;
  END A2[6]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2370 0.0010 24.4370 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2370 0.0010 24.4370 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2370 0.0000 24.4370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2370 0.0000 24.4370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2370 0.0000 24.4370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1514 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1514 LAYER M4 ;
    ANTENNAMAXAREACAR 69.5861 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1514 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1514 LAYER M5 ;
    ANTENNAMAXAREACAR 76.79102 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[15]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5540 0.0000 23.7540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5540 0.0000 23.7540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5540 0.0000 23.7540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5540 0.0000 23.7540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5540 0.0000 23.7540 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[6]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8690 0.0000 23.0690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9730 0.0000 27.1730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9730 0.0000 27.1730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9730 0.0000 27.1730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9730 0.0000 27.1730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9730 0.0000 27.1730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2900 0.0000 26.4900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2900 0.0000 26.4900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2900 0.0000 26.4900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2900 0.0000 26.4900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2900 0.0000 26.4900 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[2]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6050 0.0000 25.8050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6050 0.0000 25.8050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6050 0.0000 25.8050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6050 0.0000 25.8050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.9220 0.0000 25.1220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.9220 0.0000 25.1220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.9220 0.0000 25.1220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.9220 0.0000 25.1220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.9220 0.0000 25.1220 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[15]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6580 0.0000 27.8580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6580 0.0000 27.8580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6580 0.0000 27.8580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6580 0.0000 27.8580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6580 0.0000 27.8580 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[4]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3940 0.0000 30.5940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3940 0.0000 30.5940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3940 0.0000 30.5940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3940 0.0000 30.5940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3940 0.0000 30.5940 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7090 0.0000 29.9090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7090 0.0000 29.9090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7090 0.0000 29.9090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7090 0.0000 29.9090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7090 0.0000 29.9090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.0260 0.0000 29.2260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.0260 0.0000 29.2260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.0260 0.0000 29.2260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.0260 0.0000 29.2260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.0260 0.0000 29.2260 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
  END O2[11]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3410 0.0000 28.5410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3410 0.0000 28.5410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3410 0.0000 28.5410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3410 0.0000 28.5410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3410 0.0000 28.5410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1300 0.0000 33.3300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1300 0.0000 33.3300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1300 0.0000 33.3300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1300 0.0000 33.3300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1300 0.0000 33.3300 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4450 0.0000 32.6450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4450 0.0000 32.6450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4450 0.0000 32.6450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4450 0.0000 32.6450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4450 0.0000 32.6450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7620 0.0000 31.9620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7620 0.0000 31.9620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7620 0.0000 31.9620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7620 0.0000 31.9620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7620 0.0000 31.9620 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0770 0.0000 31.2770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0770 0.0000 31.2770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0770 0.0000 31.2770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0770 0.0000 31.2770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0770 0.0000 31.2770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8130 0.0000 34.0130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.283781 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.283781 LAYER M3 ;
    ANTENNAMAXAREACAR 62.38069 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59563 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.81008 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 125.8640 87.6300 126.0640 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 125.8640 87.6300 126.0640 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 125.8640 87.6300 126.0640 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 125.8640 87.6300 126.0640 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 125.8640 87.6300 126.0640 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2887 LAYER M1 ;
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 124.2500 87.6300 124.4500 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 124.2500 87.6300 124.4500 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 124.2500 87.6300 124.4500 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 124.2500 87.6300 124.4500 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 124.2500 87.6300 124.4500 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2887 LAYER M1 ;
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.4300 117.0440 87.6300 117.2440 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.4300 117.0440 87.6300 117.2440 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.4300 117.0440 87.6300 117.2440 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.4300 117.0440 87.6300 117.2440 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.4300 117.0440 87.6300 117.2440 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.2887 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2887 LAYER M1 ;
  END A1[3]
  OBS
    LAYER M1 ;
      RECT 0.8000 133.8920 86.8300 138.6230 ;
      RECT 0.8000 132.5320 86.8300 138.6230 ;
      RECT 0.8000 132.5320 86.8300 138.6230 ;
      RECT 0.8000 132.5320 86.8300 138.6230 ;
      RECT 0.8000 132.5320 86.8300 138.6230 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8520 ;
      RECT 0.8000 132.5320 86.8300 136.8160 ;
      RECT 0.8000 135.0620 86.8300 135.4520 ;
      RECT 0.0000 125.1140 0.8000 125.2350 ;
      RECT 0.0000 116.2820 0.8000 116.4000 ;
      RECT 21.3800 0.0000 22.2690 0.8000 ;
      RECT 86.1290 136.8520 87.6300 138.6230 ;
      RECT 86.8300 136.8160 87.6300 136.8520 ;
      RECT 0.0000 123.6500 3.0010 123.7140 ;
      RECT 0.0000 136.8520 1.5010 138.6950 ;
      RECT 0.0000 114.8320 3.0010 114.8820 ;
      RECT 0.0000 133.9320 1.5010 135.4520 ;
      RECT 0.0000 129.5310 86.8300 132.5320 ;
      RECT 86.8300 125.0500 87.6300 125.2640 ;
      RECT 86.8300 133.8920 87.6300 135.0620 ;
      RECT 86.8300 116.2320 87.6300 116.4440 ;
      RECT 0.8000 140.0230 87.6300 143.0240 ;
      RECT 0.0000 0.0000 19.9800 9.2200 ;
      RECT 0.0000 0.0000 19.9800 0.8000 ;
      RECT 0.0000 16.2280 86.8300 16.2340 ;
      RECT 0.0000 10.6210 86.8300 16.2340 ;
      RECT 0.0000 10.6210 86.8300 16.2340 ;
      RECT 0.0000 10.6210 86.8300 16.2340 ;
      RECT 0.0000 10.6210 87.6300 16.2280 ;
      RECT 0.8000 10.6200 87.6300 16.2280 ;
      RECT 0.8000 10.6200 87.6300 16.2280 ;
      RECT 0.8000 10.6200 87.6300 16.2280 ;
      RECT 0.8000 9.2210 86.8300 16.2280 ;
      RECT 0.8000 9.2210 86.8300 16.2280 ;
      RECT 0.8000 9.2210 86.8300 16.2280 ;
      RECT 0.8000 10.6200 87.6300 10.6210 ;
      RECT 0.8000 9.2210 86.8300 10.6200 ;
      RECT 0.0000 31.8380 86.8300 31.8400 ;
      RECT 0.0000 18.1680 86.8300 31.8400 ;
      RECT 0.0000 18.1680 86.8300 31.8400 ;
      RECT 0.0000 18.1680 86.8300 31.8400 ;
      RECT 0.0000 18.1680 87.6300 31.8380 ;
      RECT 0.8000 18.0900 87.6300 18.1680 ;
      RECT 0.8000 16.2340 86.8300 18.0900 ;
      RECT 0.8000 107.6040 86.8300 108.9960 ;
      RECT 0.8000 107.5960 87.6300 107.6040 ;
      RECT 0.0000 33.2400 87.6300 107.5960 ;
      RECT 0.8000 33.2400 86.8300 108.9960 ;
      RECT 0.8000 33.2400 86.8300 108.9960 ;
      RECT 0.8000 33.2400 86.8300 108.9960 ;
      RECT 0.8000 33.2400 87.6300 107.6040 ;
      RECT 0.8000 33.2400 87.6300 107.6040 ;
      RECT 0.8000 33.2400 87.6300 107.6040 ;
      RECT 0.8000 33.2380 87.6300 107.5960 ;
      RECT 0.8000 33.2380 87.6300 107.5960 ;
      RECT 0.8000 33.2380 87.6300 107.5960 ;
      RECT 0.8000 31.8400 86.8300 107.5960 ;
      RECT 0.8000 31.8400 86.8300 107.5960 ;
      RECT 0.8000 31.8400 86.8300 107.5960 ;
      RECT 0.8000 33.2380 87.6300 33.2400 ;
      RECT 0.8000 31.8400 86.8300 33.2380 ;
      RECT 0.0000 9.2200 86.8300 9.2210 ;
      RECT 0.0000 0.8000 86.8300 9.2210 ;
      RECT 0.0000 0.8000 86.8300 9.2210 ;
      RECT 0.0000 0.8000 86.8300 9.2210 ;
      RECT 0.0000 0.8000 87.6300 9.2200 ;
      RECT 67.6440 0.0000 87.6300 9.2200 ;
      RECT 67.6440 0.0000 87.6300 0.8000 ;
      RECT 0.8000 136.8520 86.8300 138.6230 ;
      RECT 0.0000 109.0040 87.6300 114.8320 ;
      RECT 0.0000 108.9960 86.8300 109.0040 ;
      RECT 0.0000 117.8000 86.8300 123.6500 ;
      RECT 0.0000 117.8440 87.6300 123.6500 ;
      RECT 0.0000 117.8000 86.8300 117.8440 ;
      RECT 0.0000 126.6350 86.8300 132.4920 ;
      RECT 0.0000 126.6640 87.6300 132.4920 ;
      RECT 0.0000 126.6350 86.8300 126.6640 ;
      RECT 0.8000 123.7140 86.8300 132.4920 ;
      RECT 0.8000 123.7140 86.8300 132.4920 ;
      RECT 0.8000 123.6500 86.8300 132.4920 ;
      RECT 0.8000 123.6500 86.8300 126.6640 ;
      RECT 0.8000 123.6500 86.8300 126.6640 ;
      RECT 0.8000 123.6500 86.8300 126.6640 ;
      RECT 0.8000 123.6500 86.8300 126.6640 ;
      RECT 0.8000 123.6500 86.8300 126.6640 ;
      RECT 0.8000 123.6500 86.8300 126.6640 ;
      RECT 0.8000 114.8820 86.8300 123.6500 ;
      RECT 0.8000 114.8820 86.8300 123.6500 ;
      RECT 0.8000 114.8320 86.8300 123.6500 ;
      RECT 0.8000 114.8320 86.8300 117.8440 ;
      RECT 0.8000 114.8320 86.8300 117.8440 ;
      RECT 0.8000 114.8320 86.8300 117.8440 ;
      RECT 0.8000 114.8320 86.8300 117.8440 ;
      RECT 0.8000 114.8320 86.8300 117.8440 ;
      RECT 0.8000 114.8320 86.8300 117.8440 ;
      RECT 0.8000 138.6230 86.8300 138.6950 ;
      RECT 0.8000 135.4520 86.8300 138.6950 ;
      RECT 0.8000 135.4520 86.8300 138.6950 ;
      RECT 0.0000 140.0950 87.6300 146.0250 ;
      RECT 0.8000 133.8920 86.8300 140.0230 ;
      RECT 0.8000 132.5320 86.8300 140.0230 ;
      RECT 0.8000 132.5320 86.8300 138.6950 ;
      RECT 0.8000 133.8920 86.8300 138.6230 ;
    LAYER PO ;
      RECT 0.0000 0.0000 87.6300 146.0250 ;
    LAYER M2 ;
      RECT 67.7440 0.0000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 0.9000 ;
      RECT 0.0000 126.7640 87.6300 132.3920 ;
      RECT 0.0000 126.7350 86.7300 126.7640 ;
      RECT 0.9000 123.6140 86.7300 126.7640 ;
      RECT 0.9000 134.9620 86.7300 135.3520 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 136.9160 ;
      RECT 0.0000 140.1950 87.6300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 136.9520 86.7300 140.1950 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 21.4800 0.0000 22.1690 0.9000 ;
      RECT 0.0000 129.4310 86.7300 132.4320 ;
      RECT 0.0000 134.0320 0.9000 135.3520 ;
      RECT 0.0000 136.9520 1.5010 138.5950 ;
      RECT 86.7300 133.9920 87.6300 134.9620 ;
      RECT 86.1290 136.9160 87.6300 138.5230 ;
      RECT 84.6290 140.1230 87.6300 140.1950 ;
      RECT 0.0000 0.0000 19.8800 9.1200 ;
      RECT 0.0000 0.0000 19.8800 0.9000 ;
      RECT 0.0000 117.9440 87.6300 123.5500 ;
      RECT 0.0000 123.5500 86.7300 123.6140 ;
      RECT 0.0000 117.9440 86.7300 123.6140 ;
      RECT 0.9000 123.6140 86.7300 126.7350 ;
      RECT 0.9000 117.9440 86.7300 126.7350 ;
      RECT 0.0000 18.2680 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 18.2680 ;
      RECT 0.9000 16.1340 86.7300 18.1900 ;
      RECT 0.0000 16.1280 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 87.6300 16.1280 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 10.7210 ;
      RECT 0.9000 9.1210 86.7300 10.7200 ;
      RECT 0.0000 117.9000 86.7300 117.9440 ;
      RECT 0.0000 114.7320 86.7300 114.7820 ;
      RECT 0.0000 109.1040 86.7300 114.7820 ;
      RECT 0.0000 109.1040 87.6300 114.7320 ;
      RECT 0.9000 114.7820 86.7300 117.9440 ;
      RECT 0.9000 114.7820 86.7300 117.9000 ;
      RECT 0.9000 109.1040 86.7300 117.9000 ;
      RECT 0.0000 109.0960 86.7300 109.1040 ;
      RECT 0.0000 31.7380 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.9000 33.3380 87.6300 33.3400 ;
      RECT 0.9000 31.7400 86.7300 33.3380 ;
      RECT 0.0000 33.3400 87.6300 107.4960 ;
      RECT 0.9000 107.5040 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 107.4960 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 31.7400 86.7300 107.4960 ;
      RECT 0.9000 31.7400 86.7300 107.4960 ;
      RECT 0.9000 31.7400 86.7300 107.4960 ;
      RECT 0.0000 9.1200 86.7300 9.1210 ;
      RECT 0.0000 0.9000 86.7300 9.1210 ;
      RECT 0.0000 0.9000 86.7300 9.1210 ;
      RECT 0.0000 0.9000 86.7300 9.1210 ;
      RECT 0.0000 0.9000 87.6300 9.1200 ;
    LAYER M3 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.9000 33.3380 87.6300 33.3400 ;
      RECT 0.9000 31.7400 86.7300 33.3380 ;
      RECT 0.0000 33.3400 87.6300 107.4960 ;
      RECT 0.9000 107.5040 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 107.4960 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 31.7400 86.7300 107.4960 ;
      RECT 0.9000 31.7400 86.7300 107.4960 ;
      RECT 0.9000 31.7400 86.7300 107.4960 ;
      RECT 0.0000 9.1200 86.7300 9.1210 ;
      RECT 0.0000 0.9000 86.7300 9.1210 ;
      RECT 0.0000 0.9000 86.7300 9.1210 ;
      RECT 0.0000 0.9000 86.7300 9.1210 ;
      RECT 0.0000 0.9000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 0.9000 ;
      RECT 0.0000 126.7640 87.6300 132.3920 ;
      RECT 0.0000 126.7350 86.7300 126.7640 ;
      RECT 0.9000 123.6140 86.7300 126.7640 ;
      RECT 0.9000 134.9620 86.7300 135.3520 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 136.9160 ;
      RECT 0.0000 140.1950 87.6300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 136.9520 86.7300 140.1950 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 21.4800 0.0000 22.1690 0.9000 ;
      RECT 0.0000 136.9520 1.5010 138.5950 ;
      RECT 0.0000 134.0320 0.9000 135.3520 ;
      RECT 0.0000 129.4310 86.7300 132.4320 ;
      RECT 84.6290 140.1230 87.6300 140.1950 ;
      RECT 86.1290 136.9160 87.6300 138.5230 ;
      RECT 86.7300 133.9920 87.6300 134.9620 ;
      RECT 0.0000 0.0000 19.8800 9.1200 ;
      RECT 0.0000 0.0000 19.8800 0.9000 ;
      RECT 0.0000 117.9440 87.6300 123.5500 ;
      RECT 0.0000 123.5500 86.7300 123.6140 ;
      RECT 0.0000 117.9440 86.7300 123.6140 ;
      RECT 0.9000 123.6140 86.7300 126.7350 ;
      RECT 0.9000 117.9440 86.7300 126.7350 ;
      RECT 0.0000 18.2680 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 18.2680 ;
      RECT 0.9000 16.1340 86.7300 18.1900 ;
      RECT 0.0000 16.1280 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 87.6300 16.1280 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 10.7210 ;
      RECT 0.9000 9.1210 86.7300 10.7200 ;
      RECT 0.0000 117.9000 86.7300 117.9440 ;
      RECT 0.0000 114.7320 86.7300 114.7820 ;
      RECT 0.0000 109.1040 86.7300 114.7820 ;
      RECT 0.0000 109.1040 87.6300 114.7320 ;
      RECT 0.9000 114.7820 86.7300 117.9440 ;
      RECT 0.9000 114.7820 86.7300 117.9000 ;
      RECT 0.9000 109.1040 86.7300 117.9000 ;
      RECT 0.0000 109.0960 86.7300 109.1040 ;
      RECT 0.0000 31.7380 86.7300 31.7400 ;
    LAYER M4 ;
      RECT 0.0000 109.0960 86.7300 109.1040 ;
      RECT 0.9000 107.5040 86.7300 109.0960 ;
      RECT 0.0000 31.7380 86.7300 31.7400 ;
      RECT 0.0000 16.1280 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 10.7210 ;
      RECT 0.0000 33.3400 87.6300 107.4960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 107.4960 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 33.3400 ;
      RECT 0.9000 31.7400 86.7300 33.3380 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 18.2680 ;
      RECT 0.9000 16.1340 86.7300 18.1900 ;
      RECT 0.0000 9.1200 86.7300 9.1210 ;
      RECT 0.0000 0.9010 86.7300 9.1210 ;
      RECT 0.0000 0.9010 86.7300 9.1210 ;
      RECT 0.0000 0.9010 86.7300 9.1210 ;
      RECT 0.0000 0.9010 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 0.9010 ;
      RECT 67.7440 0.0000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 0.9000 ;
      RECT 0.0000 126.7640 87.6300 132.3920 ;
      RECT 0.0000 126.7350 86.7300 126.7640 ;
      RECT 0.9000 123.6140 86.7300 126.7640 ;
      RECT 0.9000 134.9620 86.7300 135.3520 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 138.5230 ;
      RECT 0.9000 132.4320 86.7300 136.9160 ;
      RECT 0.0000 140.1950 87.6300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 135.3520 86.7300 146.0250 ;
      RECT 0.9000 136.9520 86.7300 140.1950 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 21.4800 0.0000 22.1690 0.9000 ;
      RECT 0.0000 136.9520 1.5010 138.5950 ;
      RECT 0.0000 134.0320 0.9000 135.3520 ;
      RECT 0.0000 129.4310 86.7300 132.4320 ;
      RECT 84.6290 140.1230 87.6300 140.1950 ;
      RECT 86.1290 136.9160 87.6300 138.5230 ;
      RECT 86.7300 133.9920 87.6300 134.9620 ;
      RECT 0.0000 0.0000 19.8800 0.9000 ;
      RECT 0.0000 0.9000 23.5370 0.9010 ;
      RECT 0.0000 0.0000 19.8800 9.1200 ;
      RECT 0.0000 0.0000 19.8800 9.1200 ;
      RECT 0.0000 0.9000 23.5370 9.1200 ;
      RECT 0.0000 0.9000 23.5370 9.1200 ;
      RECT 0.0000 0.9000 23.5370 9.1200 ;
      RECT 0.0000 117.9440 87.6300 123.5500 ;
      RECT 0.0000 109.1040 87.6300 114.7320 ;
      RECT 0.0000 117.9000 86.7300 117.9440 ;
      RECT 0.0000 114.7320 86.7300 114.7820 ;
      RECT 0.0000 109.1040 86.7300 114.7820 ;
      RECT 0.9000 114.7820 86.7300 117.9440 ;
      RECT 0.9000 114.7820 86.7300 117.9000 ;
      RECT 0.9000 109.1040 86.7300 117.9000 ;
      RECT 0.0000 123.5500 86.7300 123.6140 ;
      RECT 0.0000 117.9440 86.7300 123.6140 ;
      RECT 0.9000 123.6140 86.7300 126.7350 ;
      RECT 0.9000 117.9440 86.7300 126.7350 ;
      RECT 0.9000 9.1210 86.7300 10.7200 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 87.6300 146.0250 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 87.6300 146.0250 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 87.6300 146.0250 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 87.6300 146.0250 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 87.6300 146.0250 ;
    LAYER M5 ;
      RECT 0.0000 145.0250 0.3080 146.0250 ;
      RECT 21.4800 0.0000 22.1690 0.9000 ;
      RECT 87.0580 145.0250 87.6300 146.0250 ;
      RECT 0.0000 129.4310 86.7300 132.4320 ;
      RECT 0.0000 136.9520 1.5010 138.5950 ;
      RECT 0.0000 134.0320 0.9000 135.3520 ;
      RECT 0.9000 140.1230 87.6300 143.1240 ;
      RECT 86.1290 136.9160 87.6300 138.5230 ;
      RECT 86.7300 133.9920 87.6300 134.9620 ;
      RECT 0.0000 0.0000 19.8800 9.1200 ;
      RECT 0.0000 0.0000 19.8800 9.1200 ;
      RECT 0.0000 0.9000 23.5370 9.1200 ;
      RECT 0.0000 0.9000 23.5370 9.1200 ;
      RECT 0.0000 0.9000 23.5370 9.1200 ;
      RECT 0.0000 0.9000 23.5370 0.9010 ;
      RECT 0.0000 0.0000 19.8800 0.9000 ;
      RECT 0.0000 117.9440 87.6300 123.5500 ;
      RECT 0.0000 109.1040 87.6300 114.7320 ;
      RECT 0.0000 117.9000 86.7300 117.9440 ;
      RECT 0.0000 114.7320 86.7300 114.7820 ;
      RECT 0.0000 109.1040 86.7300 114.7820 ;
      RECT 0.9000 114.7820 86.7300 117.9440 ;
      RECT 0.9000 114.7820 86.7300 117.9000 ;
      RECT 0.9000 109.1040 86.7300 117.9000 ;
      RECT 0.0000 123.5500 86.7300 123.6140 ;
      RECT 0.0000 117.9440 86.7300 123.6140 ;
      RECT 0.9000 123.6140 86.7300 126.7350 ;
      RECT 0.9000 117.9440 86.7300 126.7350 ;
      RECT 0.9000 9.1210 86.7300 10.7200 ;
      RECT 0.0000 109.0960 86.7300 109.1040 ;
      RECT 0.9000 107.5040 86.7300 109.0960 ;
      RECT 0.0000 31.7380 86.7300 31.7400 ;
      RECT 0.0000 16.1280 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 86.7300 16.1340 ;
      RECT 0.0000 10.7210 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 9.1210 86.7300 16.1280 ;
      RECT 0.9000 10.7200 87.6300 10.7210 ;
      RECT 0.0000 33.3400 87.6300 107.4960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 33.3400 86.7300 109.0960 ;
      RECT 0.9000 107.4960 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3400 87.6300 107.5040 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 107.4960 ;
      RECT 0.9000 33.3380 87.6300 33.3400 ;
      RECT 0.9000 31.7400 86.7300 33.3380 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 86.7300 31.7400 ;
      RECT 0.0000 18.2680 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 10.7210 86.7300 31.7380 ;
      RECT 0.9000 18.1900 87.6300 18.2680 ;
      RECT 0.9000 16.1340 86.7300 18.1900 ;
      RECT 0.0000 9.1200 86.7300 9.1210 ;
      RECT 0.0000 0.9010 86.7300 9.1210 ;
      RECT 0.0000 0.9010 86.7300 9.1210 ;
      RECT 0.0000 0.9010 86.7300 9.1210 ;
      RECT 0.0000 0.9010 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 9.1200 ;
      RECT 25.1370 0.9000 87.6300 0.9010 ;
      RECT 67.7440 0.0000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 9.1200 ;
      RECT 67.7440 0.0000 87.6300 0.9000 ;
      RECT 0.9000 134.9620 86.7300 135.3520 ;
      RECT 0.9000 138.5230 86.7300 138.5950 ;
      RECT 0.9000 135.3520 86.7300 138.5950 ;
      RECT 0.9000 135.3520 86.7300 138.5950 ;
      RECT 0.9000 135.3520 86.7300 138.5950 ;
      RECT 0.0000 140.1950 87.6300 145.0250 ;
      RECT 0.9000 136.9160 86.7300 140.1230 ;
      RECT 0.9000 136.9160 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.9000 135.3520 86.7300 140.1230 ;
      RECT 0.0000 126.7640 87.6300 132.3920 ;
      RECT 0.0000 126.7350 86.7300 126.7640 ;
      RECT 0.9000 132.4320 86.7300 136.9160 ;
      RECT 0.9000 123.6140 86.7300 126.7640 ;
  END
END SRAMLP2RW128x16

MACRO SRAMLP2RW128x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 131.406 BY 154.678 ;
  SYMMETRY X Y R90 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 129.7090 154.3780 130.0080 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.8100 154.3780 129.1100 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.4090 154.3780 15.7090 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.9080 154.3780 11.2090 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.8080 154.3780 12.1090 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.0080 154.3780 1.3080 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9090 154.3780 2.2080 154.6780 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.1580 154.3780 4.4590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2580 154.3780 3.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3590 154.3780 2.6590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4580 154.3780 1.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0580 154.3780 5.3590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5580 154.3780 9.8590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6580 154.3780 8.9590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7590 154.3780 8.0580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8590 154.3780 7.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9590 154.3780 6.2590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3590 154.3780 11.6580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4590 154.3780 10.7590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0580 154.3780 14.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1590 154.3780 13.4590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2580 154.3780 12.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5580 154.3780 18.8590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6580 154.3780 17.9590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7580 154.3780 17.0590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8580 154.3780 16.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9590 154.3780 15.2580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2580 154.3780 21.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3590 154.3780 20.6590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1580 154.3780 22.4590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9590 154.3780 24.2580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0590 154.3780 23.3590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4590 154.3780 19.7590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7580 154.3780 26.0580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6590 154.3780 26.9590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5580 154.3780 27.8580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4590 154.3780 28.7590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8580 154.3780 25.1590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9590 154.3780 33.2590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1580 154.3780 31.4590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3590 154.3780 29.6580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2590 154.3780 30.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0580 154.3780 32.3590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8590 154.3780 34.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4580 154.3780 37.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6580 154.3780 35.9590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5580 154.3780 36.8590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3580 154.3780 38.6580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7590 154.3780 35.0580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8580 154.3780 43.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2590 154.3780 39.5590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1580 154.3780 40.4570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9580 154.3780 42.2580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0590 154.3780 41.3600 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3580 154.3780 47.6580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2590 154.3780 48.5590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4580 154.3780 46.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7590 154.3780 44.0590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5590 154.3780 45.8600 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6580 154.3780 44.9570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8580 154.3780 52.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1580 154.3780 49.4570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0590 154.3780 50.3600 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7590 154.3780 53.0590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9580 154.3780 51.2580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2580 154.3780 57.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4580 154.3780 55.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5580 154.3780 54.8580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6580 154.3780 53.9580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3590 154.3780 56.6590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6570 154.3780 62.9570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7580 154.3780 62.0580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8580 154.3780 61.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0580 154.3780 59.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1580 154.3780 58.4580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9590 154.3780 60.2590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1570 154.3780 67.4570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2580 154.3780 66.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3570 154.3780 65.6570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4570 154.3780 64.7570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5580 154.3780 63.8580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6580 154.3780 71.9580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7590 154.3780 71.0590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8570 154.3780 70.1570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9570 154.3780 69.2570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0580 154.3780 68.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1570 154.3780 76.4570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2580 154.3780 75.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3580 154.3780 74.6580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4580 154.3780 73.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.0580 154.3780 77.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5590 154.3780 72.8590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6580 154.3780 80.9580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7600 154.3780 80.0600 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8570 154.3780 79.1570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9570 154.3780 78.2570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5590 154.3780 81.8590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.9570 154.3780 87.2570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1570 154.3780 85.4570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2580 154.3780 84.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3580 154.3780 83.6580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4580 154.3780 82.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0580 154.3780 86.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.4580 154.3780 91.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.5580 154.3780 90.8580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.6580 154.3780 89.9580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.8580 154.3780 88.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.7590 154.3780 89.0590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.0580 154.3780 95.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.1570 154.3780 94.4570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.3570 154.3780 92.6570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.9590 154.3780 96.2590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.2580 154.3780 93.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.3570 154.3780 101.6570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.5570 154.3780 99.8570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.6580 154.3780 98.9580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.7580 154.3780 98.0580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.8580 154.3780 97.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.4580 154.3780 100.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.8590 154.3780 106.1590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.9590 154.3780 105.2590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.0590 154.3780 104.3590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.2590 154.3780 102.5590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.1600 154.3780 103.4600 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.4580 154.3780 109.7580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.5580 154.3780 108.8580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.7580 154.3780 107.0580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.3590 154.3780 110.6590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.6590 154.3780 107.9590 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.7570 154.3780 116.0570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.9570 154.3780 114.2570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.0580 154.3780 113.3580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.1580 154.3780 112.4580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.2580 154.3780 111.5580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.8580 154.3780 115.1580 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.2560 154.3780 120.5560 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.3560 154.3780 119.6560 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.4560 154.3780 118.7560 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.6560 154.3780 116.9560 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.5570 154.3780 117.8570 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.7550 154.3780 125.0550 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.0560 154.3780 122.3560 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.8540 154.3780 124.1540 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.9550 154.3780 123.2550 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.6540 154.3780 125.9540 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.5540 154.3780 126.8540 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.4540 154.3780 127.7540 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.3530 154.3780 128.6530 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.1530 154.3780 130.4530 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.2540 154.3780 129.5540 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.1550 154.3780 121.4550 154.6780 ;
    END
  END VSS

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.9600 0.0020 91.1600 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.9600 0.0020 91.1600 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.9600 0.0020 91.1600 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.9600 0.0020 91.1600 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.9600 0.0020 91.1600 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[29]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.5920 0.0020 89.7920 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.5920 0.0020 89.7920 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.5920 0.0020 89.7920 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.5920 0.0020 89.7920 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.5920 0.0020 89.7920 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[22]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.2240 0.0020 88.4240 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.2240 0.0020 88.4240 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.2240 0.0020 88.4240 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.2240 0.0020 88.4240 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.2240 0.0020 88.4240 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[26]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.3020 0.0000 90.5020 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[29]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.9340 0.0000 89.1340 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[22]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6960 0.0020 93.8960 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6960 0.0020 93.8960 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6960 0.0020 93.8960 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6960 0.0020 93.8960 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6960 0.0020 93.8960 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[15]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.3280 0.0020 92.5280 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.3280 0.0020 92.5280 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.3280 0.0020 92.5280 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.3280 0.0020 92.5280 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.3280 0.0020 92.5280 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[21]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.4060 0.0000 94.6060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[27]

  PIN DS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 144.7800 0.2000 144.9800 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 144.7800 0.2000 144.9800 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 144.7800 0.2000 144.9800 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 144.7800 0.2000 144.9800 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 144.7800 0.2000 144.9800 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAGATEAREA 0.2256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.381834 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.381834 LAYER M2 ;
    ANTENNAMAXAREACAR 6.258323 LAYER M2 ;
    ANTENNAGATEAREA 0.8058 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 16.78506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.78506 LAYER M3 ;
    ANTENNAMAXAREACAR 32.34911 LAYER M3 ;
    ANTENNAGATEAREA 0.8058 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 42.3474 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.3474 LAYER M4 ;
    ANTENNAMAXAREACAR 84.90234 LAYER M4 ;
    ANTENNAGATEAREA 54.1422 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 11289.29 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 11289.29 LAYER M5 ;
    ANTENNAMAXAREACAR 291.9471 LAYER M5 ;
    ANTENNAGATEAREA 54.1422 LAYER M6 ;
    ANTENNAGATEAREA 54.1422 LAYER M7 ;
    ANTENNAGATEAREA 54.1422 LAYER M8 ;
    ANTENNAGATEAREA 54.1422 LAYER M9 ;
    ANTENNAGATEAREA 54.1422 LAYER MRDL ;
  END DS2

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.6700 0.0000 91.8700 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[21]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.7740 0.0000 95.9740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[20]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.8010 0.0020 98.0010 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.8010 0.0020 98.0010 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.8010 0.0020 98.0010 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.8010 0.0020 98.0010 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.8010 0.0020 98.0010 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[24]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.4320 0.0020 96.6320 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.4320 0.0020 96.6320 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.4320 0.0020 96.6320 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.4320 0.0020 96.6320 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.4320 0.0020 96.6320 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[20]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.1420 0.0000 97.3420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[24]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.0640 0.0020 95.2640 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.0640 0.0020 95.2640 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.0640 0.0020 95.2640 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.0640 0.0020 95.2640 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.0640 0.0020 95.2640 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[27]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.5180 0.0000 72.7180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[30]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.1500 0.0000 71.3500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[19]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.9120 0.0020 76.1120 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[13]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.2540 0.0000 75.4540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[13]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.5440 0.0020 74.7440 0.2020 ;
    END
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[5]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.2800 0.0020 77.4800 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[1]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.6220 0.0000 76.8220 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[1]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.3840 0.0020 81.5840 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.0160 0.0020 80.2160 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[11]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.6480 0.0020 78.8480 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[28]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.7820 0.0000 69.9820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[14]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.3580 0.0000 79.5580 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[11]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.9900 0.0000 78.1900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[28]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.0940 0.0000 82.2940 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[25]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.1980 0.0000 86.3980 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[31]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.8300 0.0000 85.0300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.8300 0.0000 85.0300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.8300 0.0000 85.0300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.8300 0.0000 85.0300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.8300 0.0000 85.0300 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[0]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.4620 0.0000 83.6620 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[23]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.8560 0.0020 87.0560 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.8560 0.0020 87.0560 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.8560 0.0020 87.0560 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.8560 0.0020 87.0560 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.8560 0.0020 87.0560 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[31]

  PIN O2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0940 0.0020 59.2940 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0940 0.0020 59.2940 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0940 0.0020 59.2940 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0940 0.0020 59.2940 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0940 0.0020 59.2940 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[10]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1720 0.0000 61.3720 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[3]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.8040 0.0000 60.0040 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.4360 0.0000 58.6360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[10]

  PIN O2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.7260 0.0020 57.9260 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.7260 0.0020 57.9260 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.7260 0.0020 57.9260 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.7260 0.0020 57.9260 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.7260 0.0020 57.9260 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[17]

  PIN O2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1980 0.0020 63.3980 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1980 0.0020 63.3980 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1980 0.0020 63.3980 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1980 0.0020 63.3980 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1980 0.0020 63.3980 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[16]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.5400 0.0000 62.7400 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[16]

  PIN O2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.9340 0.0020 66.1340 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.9340 0.0020 66.1340 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.9340 0.0020 66.1340 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.9340 0.0020 66.1340 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.9340 0.0020 66.1340 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[12]

  PIN O2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5660 0.0020 64.7660 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5660 0.0020 64.7660 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5660 0.0020 64.7660 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5660 0.0020 64.7660 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5660 0.0020 64.7660 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[8]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2760 0.0000 65.4760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[12]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.9080 0.0000 64.1080 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[8]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.0720 0.0020 69.2720 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[6]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.7040 0.0020 67.9040 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[2]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.0460 0.0000 67.2460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[2]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.4140 0.0000 68.6140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[6]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.4400 0.0020 70.6400 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[14]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.1760 0.0020 73.3760 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[30]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.8080 0.0020 72.0080 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[19]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.8860 0.0000 74.0860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[5]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 141.8340 131.4060 142.0340 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 141.8340 131.4060 142.0340 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 141.8340 131.4060 142.0340 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 141.8340 131.4060 142.0340 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 141.8340 131.4060 142.0340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.28814 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28814 LAYER M1 ;
  END A1[0]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 9.8960 0.2000 10.0960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15256 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15256 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56742 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56742 LAYER M2 ;
    ANTENNAMAXAREACAR 11.76674 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.80361 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.84041 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.87714 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 16.9090 0.2000 17.1090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.40684 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40684 LAYER M4 ;
    ANTENNAMAXAREACAR 13.56469 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.70587 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB2

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 17.4430 0.2000 17.6430 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15736 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0894 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30916 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30916 LAYER M4 ;
    ANTENNAMAXAREACAR 6.377295 LAYER M4 ;
    ANTENNAGATEAREA 0.0894 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 8.072623 LAYER M5 ;
    ANTENNAGATEAREA 0.0894 LAYER M6 ;
    ANTENNAGATEAREA 0.0894 LAYER M7 ;
    ANTENNAGATEAREA 0.0894 LAYER M8 ;
    ANTENNAGATEAREA 0.0894 LAYER M9 ;
    ANTENNAGATEAREA 0.0894 LAYER MRDL ;
  END CE2

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 41.1530 0.2000 41.3530 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 41.1530 0.2000 41.3530 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 41.1530 0.2000 41.3530 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 41.1530 0.2000 41.3530 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 41.1530 0.2000 41.3530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.296184 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296184 LAYER M1 ;
    ANTENNAGATEAREA 0.021 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.84244 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.84244 LAYER M2 ;
    ANTENNAMAXAREACAR 47.09487 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 54.31081 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 61.52628 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 68.74126 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A2[6]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 124.2060 0.2000 124.4060 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 124.2060 0.2000 124.4060 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 124.2060 0.2000 124.4060 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 124.2060 0.2000 124.4060 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 124.2060 0.2000 124.4060 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288456 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288456 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72196 LAYER M2 ;
    ANTENNAMAXAREACAR 21.1402 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.28088 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.42129 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.56142 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[4]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 125.7240 0.2000 125.9240 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 125.7240 0.2000 125.9240 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 125.7240 0.2000 125.9240 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 125.7240 0.2000 125.9240 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 125.7240 0.2000 125.9240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288456 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288456 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72196 LAYER M2 ;
    ANTENNAMAXAREACAR 21.13681 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.27749 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.4179 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.55804 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[3]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 133.0380 0.2000 133.2380 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 133.0380 0.2000 133.2380 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 133.0380 0.2000 133.2380 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 133.0380 0.2000 133.2380 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 133.0380 0.2000 133.2380 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288456 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288456 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72196 LAYER M2 ;
    ANTENNAMAXAREACAR 21.16053 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.30121 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.44161 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.58175 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[2]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 141.8560 0.2000 142.0560 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 141.8560 0.2000 142.0560 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 141.8560 0.2000 142.0560 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 141.8560 0.2000 142.0560 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 141.8560 0.2000 142.0560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288456 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288456 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72196 LAYER M2 ;
    ANTENNAMAXAREACAR 21.15714 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.29782 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.43823 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.57836 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 134.5590 0.2000 134.7590 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 134.5590 0.2000 134.7590 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 134.5590 0.2000 134.7590 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 134.5590 0.2000 134.7590 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 134.5590 0.2000 134.7590 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288456 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288456 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72196 LAYER M2 ;
    ANTENNAMAXAREACAR 21.1114 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.25208 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.3925 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.53263 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[1]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 41.1680 131.4060 41.3680 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 41.1680 131.4060 41.3680 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 41.1680 131.4060 41.3680 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 41.1680 131.4060 41.3680 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 41.1680 131.4060 41.3680 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15514 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.23446 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23446 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.90322 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.90322 LAYER M3 ;
    ANTENNAMAXAREACAR 51.00689 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 58.22258 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 65.43778 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END A1[6]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 116.9130 0.2000 117.1130 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 116.9130 0.2000 117.1130 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 116.9130 0.2000 117.1130 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 116.9130 0.2000 117.1130 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 116.9130 0.2000 117.1130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.288456 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.288456 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.72196 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.72196 LAYER M2 ;
    ANTENNAMAXAREACAR 21.12156 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 25.26225 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 29.40266 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.54279 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A2[5]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.3320 0.0000 54.5320 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[7]

  PIN O2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3580 0.0020 56.5580 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3580 0.0020 56.5580 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3580 0.0020 56.5580 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3580 0.0020 56.5580 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3580 0.0020 56.5580 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[18]

  PIN O2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9900 0.0020 55.1900 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9900 0.0020 55.1900 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9900 0.0020 55.1900 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9900 0.0020 55.1900 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9900 0.0020 55.1900 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[7]

  PIN O2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.6220 0.0020 53.8220 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.6220 0.0020 53.8220 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.6220 0.0020 53.8220 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.6220 0.0020 53.8220 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.6220 0.0020 53.8220 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[24]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0680 0.0000 57.2680 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[17]

  PIN O2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.8300 0.0020 62.0300 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.8300 0.0020 62.0300 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.8300 0.0020 62.0300 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.8300 0.0020 62.0300 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.8300 0.0020 62.0300 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[3]

  PIN O2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4620 0.0020 60.6620 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4620 0.0020 60.6620 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4620 0.0020 60.6620 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4620 0.0020 60.6620 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4620 0.0020 60.6620 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[9]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 124.1850 131.4060 124.3850 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 124.1850 131.4060 124.3850 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 124.1850 131.4060 124.3850 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 124.1850 131.4060 124.3850 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 124.1850 131.4060 124.3850 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.28814 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28814 LAYER M1 ;
  END A1[4]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 125.7070 131.4060 125.9070 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 125.7070 131.4060 125.9070 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 125.7070 131.4060 125.9070 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 125.7070 131.4060 125.9070 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 125.7070 131.4060 125.9070 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.28814 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28814 LAYER M1 ;
  END A1[3]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 133.0080 131.4060 133.2080 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 133.0080 131.4060 133.2080 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 133.0080 131.4060 133.2080 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 133.0080 131.4060 133.2080 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 133.0080 131.4060 133.2080 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.28814 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28814 LAYER M1 ;
  END A1[2]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 134.5340 131.4060 134.7340 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 134.5340 131.4060 134.7340 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 134.5340 131.4060 134.7340 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 134.5340 131.4060 134.7340 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 134.5340 131.4060 134.7340 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.28814 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28814 LAYER M1 ;
  END A1[1]

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 17.3650 131.4060 17.5650 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 17.3650 131.4060 17.5650 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 17.3650 131.4060 17.5650 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 17.3650 131.4060 17.5650 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 17.3650 131.4060 17.5650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.29968 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.29968 LAYER M4 ;
    ANTENNAMAXAREACAR 13.19096 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 17.62284 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE1

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 116.9040 131.4060 117.1040 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 116.9040 131.4060 117.1040 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 116.9040 131.4060 117.1040 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 116.9040 131.4060 117.1040 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 116.9040 131.4060 117.1040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.28814 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28814 LAYER M1 ;
    ANTENNAGATEAREA 21.8796 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 59.44209 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.44209 LAYER M2 ;
    ANTENNAMAXAREACAR 15.73504 LAYER M2 ;
    ANTENNAGATEAREA 23.0712 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 13.43644 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.43644 LAYER M3 ;
    ANTENNAMAXAREACAR 6.301872 LAYER M3 ;
    ANTENNAGATEAREA 23.0712 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 52.9392 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 52.9392 LAYER M4 ;
    ANTENNAMAXAREACAR 18.61201 LAYER M4 ;
    ANTENNAGATEAREA 23.0712 LAYER M5 ;
    ANTENNAGATEAREA 23.0712 LAYER M6 ;
    ANTENNAGATEAREA 23.0712 LAYER M7 ;
    ANTENNAGATEAREA 23.0712 LAYER M8 ;
    ANTENNAGATEAREA 23.0712 LAYER M9 ;
    ANTENNAGATEAREA 23.0712 LAYER MRDL ;
  END A1[5]

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 16.9030 131.4060 17.1030 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 16.9030 131.4060 17.1030 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 16.9030 131.4060 17.1030 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 16.9030 131.4060 17.1030 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 16.9030 131.4060 17.1030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.424789 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.424789 LAYER M4 ;
    ANTENNAMAXAREACAR 14.05956 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.20071 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB1

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.3760 0.0020 107.5760 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.3760 0.0020 107.5760 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[16]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 103.2720 0.0020 103.4720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.2720 0.0020 103.4720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.2720 0.0020 103.4720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.2720 0.0020 103.4720 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[10]

  PIN O2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.5180 0.0020 49.7180 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[15]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.2280 0.0000 50.4280 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[27]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8600 0.0000 49.0600 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[15]

  PIN O2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2540 0.0020 52.4540 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2540 0.0020 52.4540 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2540 0.0020 52.4540 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2540 0.0020 52.4540 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2540 0.0020 52.4540 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[20]

  PIN O2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8860 0.0020 51.0860 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[27]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9640 0.0000 53.1640 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[24]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5960 0.0000 51.7960 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[20]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.7000 0.0000 55.9000 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[18]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.0380 0.0000 93.2380 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[15]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0760 0.0020 31.2760 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[13]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.7260 0.0000 80.9260 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[4]

  PIN DS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 144.8050 131.4060 145.0050 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 144.8050 131.4060 145.0050 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 144.8050 131.4060 145.0050 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 144.8050 131.4060 145.0050 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 144.8050 131.4060 145.0050 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END DS1

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 144.4510 131.4060 144.6510 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 144.4510 131.4060 144.6510 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 144.4510 131.4060 144.6510 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 144.4510 131.4060 144.6510 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 144.4510 131.4060 144.6510 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15448 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15448 LAYER M2 ;
  END SD

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 9.8950 131.4060 10.0950 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 9.8950 131.4060 10.0950 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 9.8950 131.4060 10.0950 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 9.8950 131.4060 10.0950 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 9.8950 131.4060 10.0950 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15724 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15724 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56742 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56742 LAYER M2 ;
    ANTENNAMAXAREACAR 11.76674 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.80361 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.84041 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.87714 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB1

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 16.3090 154.3780 16.6090 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.2040 154.3780 125.5030 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.1100 154.3780 126.4090 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.5090 154.3780 5.8080 154.6780 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.6090 154.3780 4.9080 154.6780 ;
    END
    ANTENNADIFFAREA 10.5678 LAYER M5 ;
    ANTENNADIFFAREA 10.5678 LAYER M6 ;
    ANTENNADIFFAREA 10.5678 LAYER M7 ;
    ANTENNADIFFAREA 10.5678 LAYER M8 ;
    ANTENNADIFFAREA 10.5678 LAYER M9 ;
    ANTENNADIFFAREA 10.5678 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 276.3375 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 276.3375 LAYER M5 ;
  END VDDL

  PIN OEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.5780 0.0000 20.7780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.5178 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.876314 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.876314 LAYER M2 ;
    ANTENNAMAXAREACAR 6.520897 LAYER M2 ;
    ANTENNAGATEAREA 0.5178 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 6.813244 LAYER M3 ;
    ANTENNAGATEAREA 0.5178 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.105571 LAYER M4 ;
    ANTENNAGATEAREA 0.5178 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.39788 LAYER M5 ;
    ANTENNAGATEAREA 0.5178 LAYER M6 ;
    ANTENNAGATEAREA 0.5178 LAYER M7 ;
    ANTENNAGATEAREA 0.5178 LAYER M8 ;
    ANTENNAGATEAREA 0.5178 LAYER M9 ;
    ANTENNAGATEAREA 0.5178 LAYER MRDL ;
  END OEB2

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.6180 0.0000 110.8180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAGATEAREA 0.5178 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.882134 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.882134 LAYER M2 ;
    ANTENNAMAXAREACAR 6.532137 LAYER M2 ;
    ANTENNAGATEAREA 0.5178 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 6.824483 LAYER M3 ;
    ANTENNAGATEAREA 0.5178 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 7.11681 LAYER M4 ;
    ANTENNAGATEAREA 0.5178 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 7.409118 LAYER M5 ;
    ANTENNAGATEAREA 0.5178 LAYER M6 ;
    ANTENNAGATEAREA 0.5178 LAYER M7 ;
    ANTENNAGATEAREA 0.5178 LAYER M8 ;
    ANTENNAGATEAREA 0.5178 LAYER M9 ;
    ANTENNAGATEAREA 0.5178 LAYER MRDL ;
  END OEB1

  PIN LS1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.2060 147.9320 131.4060 148.1320 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.2060 147.9320 131.4060 148.1320 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.2060 147.9320 131.4060 148.1320 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.2060 147.9320 131.4060 148.1320 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.2060 147.9320 131.4060 148.1320 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.220445 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.220445 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.97624 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.01857 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.0607 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS1

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9160 0.0000 38.1160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[25]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5480 0.0000 36.7480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[4]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1800 0.0000 35.3800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[11]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8120 0.0020 34.0120 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[28]

  PIN O2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6780 0.0020 42.8780 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[31]

  PIN O2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.3100 0.0020 41.5100 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[0]

  PIN O2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9420 0.0020 40.1420 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[23]

  PIN O2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5740 0.0020 38.7740 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3880 0.0000 43.5880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[26]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0200 0.0000 42.2200 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[31]

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6520 0.0000 40.8520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[0]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2840 0.0000 39.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[23]

  PIN O2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0460 0.0020 44.2460 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[26]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4920 0.0000 47.6920 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7560 0.0000 44.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[22]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.1240 0.0000 46.3240 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[29]

  PIN O2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1500 0.0020 48.3500 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[21]

  PIN O2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7830 0.0020 46.9830 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[29]

  PIN O2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.4140 0.0020 45.6140 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[22]

  PIN O2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6300 0.0020 27.8300 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[19]

  PIN O2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2630 0.0020 26.4630 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[14]

  PIN O2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8940 0.0020 25.0940 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[6]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9720 0.0020 27.1720 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[19]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6040 0.0020 25.8040 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[14]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2360 0.0020 24.4360 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[6]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8680 0.0020 23.0680 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[2]

  PIN O2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7340 0.0020 31.9340 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[13]

  PIN O2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3660 0.0020 30.5660 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[5]

  PIN O2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9980 0.0020 29.1980 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[30]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4440 0.0020 32.6440 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[1]

  PIN LS2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 148.0090 0.2000 148.2090 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.0000 148.0090 0.2000 148.2090 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.0000 148.0090 0.2000 148.2090 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 148.0090 0.2000 148.2090 ;
    END
    PORT
      LAYER M1 ;
        RECT 0.0000 148.0090 0.2000 148.2090 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.220395 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.220395 LAYER M1 ;
    ANTENNAGATEAREA 0.0498 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.941752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.941752 LAYER M2 ;
    ANTENNAMAXAREACAR 20.8743 LAYER M2 ;
    ANTENNAGATEAREA 0.0498 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 27.97487 LAYER M3 ;
    ANTENNAGATEAREA 0.0498 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 31.0172 LAYER M4 ;
    ANTENNAGATEAREA 0.0498 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 34.05933 LAYER M5 ;
    ANTENNAGATEAREA 0.0498 LAYER M6 ;
    ANTENNAGATEAREA 0.0498 LAYER M7 ;
    ANTENNAGATEAREA 0.0498 LAYER M8 ;
    ANTENNAGATEAREA 0.0498 LAYER M9 ;
    ANTENNAGATEAREA 0.0498 LAYER MRDL ;
  END LS2

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7080 0.0020 29.9080 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[5]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3400 0.0020 28.5400 0.2020 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I2[30]

  PIN O2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 0.0020 33.3020 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[1]

  PIN O2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.2050 0.0020 37.4050 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[4]

  PIN O2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8380 0.0020 36.0380 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[11]

  PIN O2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4700 0.0020 34.6700 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[28]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.5360 0.0020 100.7360 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.5360 0.0020 100.7360 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.5360 0.0020 100.7360 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.5360 0.0020 100.7360 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.5360 0.0020 100.7360 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[18]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.1680 0.0020 99.3680 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.1680 0.0020 99.3680 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.1680 0.0020 99.3680 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.1680 0.0020 99.3680 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.1680 0.0020 99.3680 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[7]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.2460 0.0000 101.4460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.8780 0.0000 100.0780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[18]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.5100 0.0000 98.7100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[7]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.6140 0.0000 102.8140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[10]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.9820 0.0000 104.1820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[9]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.9040 0.0020 102.1040 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.9040 0.0020 102.1040 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.9040 0.0020 102.1040 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.9040 0.0020 102.1040 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.9040 0.0020 102.1040 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[17]

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.0080 0.0020 106.2080 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.0080 0.0020 106.2080 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.0080 0.0020 106.2080 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.0080 0.0020 106.2080 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.0080 0.0020 106.2080 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[3]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.6400 0.0020 104.8400 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.6400 0.0020 104.8400 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.6400 0.0020 104.8400 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.6400 0.0020 104.8400 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.6400 0.0020 104.8400 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[9]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.3500 0.0000 105.5500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[3]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.1120 0.0020 110.3120 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.1120 0.0020 110.3120 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.1120 0.0020 110.3120 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.1120 0.0020 110.3120 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.1120 0.0020 110.3120 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[12]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.7440 0.0020 108.9440 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.7440 0.0020 108.9440 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.7440 0.0020 108.9440 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.7440 0.0020 108.9440 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.7440 0.0020 108.9440 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[8]

  PIN O2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.2720 0.0020 103.4720 0.2020 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.3760 0.0020 107.5760 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.3760 0.0020 107.5760 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.3760 0.0020 107.5760 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.5220 0.0020 23.7220 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O2[2]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.0860 0.0000 108.2860 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[8]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.7180 0.0000 106.9180 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[16]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.4540 0.0000 109.6540 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28824 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28824 LAYER M3 ;
    ANTENNAMAXAREACAR 62.59302 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80795 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.02238 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[12]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.4880 0.0020 85.6880 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.4880 0.0020 85.6880 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.4880 0.0020 85.6880 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.4880 0.0020 85.6880 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.4880 0.0020 85.6880 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[0]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.1200 0.0020 84.3200 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.1200 0.0020 84.3200 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.1200 0.0020 84.3200 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.1200 0.0020 84.3200 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.1200 0.0020 84.3200 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[23]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.5360 0.0000 87.7360 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.29343 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29343 LAYER M3 ;
    ANTENNAMAXAREACAR 62.84016 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 70.05507 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.26949 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.7520 0.0020 82.9520 0.2020 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15502 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O1[25]
  OBS
    LAYER M1 ;
      RECT 0.8000 0.8020 130.6060 16.3030 ;
      RECT 0.8000 0.8020 130.6060 16.3030 ;
      RECT 0.8000 0.8020 130.6060 16.3030 ;
      RECT 110.9120 0.8000 131.4060 9.2950 ;
      RECT 110.9120 0.8000 131.4060 9.2950 ;
      RECT 110.9120 0.8000 131.4060 0.8020 ;
      RECT 111.4180 0.0000 131.4060 9.2950 ;
      RECT 111.4180 0.0000 131.4060 9.2950 ;
      RECT 111.4180 0.0000 131.4060 0.8000 ;
      RECT 0.8000 125.1070 130.6060 125.1240 ;
      RECT 0.0000 117.7130 131.4060 123.5850 ;
      RECT 0.8000 124.9850 130.6060 125.0060 ;
      RECT 0.8000 117.7040 131.4060 123.5850 ;
      RECT 0.8000 117.7040 131.4060 123.5850 ;
      RECT 0.8000 117.7040 131.4060 123.5850 ;
      RECT 0.8000 117.7040 131.4060 117.7130 ;
      RECT 0.0000 126.5240 131.4060 132.4080 ;
      RECT 0.8000 133.8080 130.6060 133.8380 ;
      RECT 0.8000 147.3320 130.6060 147.4090 ;
      RECT 0.8000 144.1800 130.6060 147.4090 ;
      RECT 0.8000 144.1800 130.6060 147.4090 ;
      RECT 0.8000 144.1800 130.6060 147.4090 ;
      RECT 0.0000 148.8090 131.4060 154.6780 ;
      RECT 0.8000 145.5800 130.6060 148.7320 ;
      RECT 0.8000 145.5800 130.6060 148.7320 ;
      RECT 0.8000 144.1800 130.6060 148.7320 ;
      RECT 0.8000 144.1800 130.6060 148.7320 ;
      RECT 0.8000 141.2560 130.6060 145.5800 ;
      RECT 0.0000 135.3590 131.4060 141.2340 ;
      RECT 66.7340 0.8000 67.1040 0.8020 ;
      RECT 0.0000 138.3350 130.6060 141.2560 ;
      RECT 0.0000 138.2550 131.4060 138.3350 ;
      RECT 0.0000 125.1070 130.6060 125.1240 ;
      RECT 0.0000 133.9340 130.6060 133.9590 ;
      RECT 0.0000 133.8380 131.4060 133.9340 ;
      RECT 0.0000 129.4370 131.4060 129.5080 ;
      RECT 0.0000 125.0060 131.4060 125.1070 ;
      RECT 0.0000 129.5080 130.6060 132.4380 ;
      RECT 0.0000 145.5800 1.5010 147.4090 ;
      RECT 0.0000 120.6050 130.6060 123.6060 ;
      RECT 0.0000 142.7350 1.5010 144.1800 ;
      RECT 0.0000 142.6560 131.4060 142.7350 ;
      RECT 0.8000 124.9850 131.4060 125.0060 ;
      RECT 0.8000 126.5070 131.4060 129.4370 ;
      RECT 0.8000 123.6060 130.6060 124.9850 ;
      RECT 0.8000 125.1240 130.6060 126.5070 ;
      RECT 0.8000 148.7320 131.4060 151.7330 ;
      RECT 0.8000 141.2560 130.6060 142.6340 ;
      RECT 0.8000 142.6340 131.4060 142.6560 ;
      RECT 0.8000 135.3340 131.4060 138.2550 ;
      RECT 0.8000 132.4380 130.6060 133.8080 ;
      RECT 0.8000 133.8080 131.4060 133.8380 ;
      RECT 0.8000 133.9590 130.6060 135.3340 ;
      RECT 21.3780 0.0000 22.2680 0.8000 ;
      RECT 66.7340 0.8000 67.1040 1.1010 ;
      RECT 129.9050 145.6050 131.4060 147.3320 ;
      RECT 130.6060 142.7350 131.4060 143.8510 ;
      RECT 0.0000 0.0000 19.9780 0.8000 ;
      RECT 0.8000 125.0060 130.6060 125.1070 ;
      RECT 0.0000 16.3030 130.6060 16.3090 ;
      RECT 0.0000 10.6960 130.6060 16.3090 ;
      RECT 0.0000 10.6960 130.6060 16.3090 ;
      RECT 0.0000 10.6960 130.6060 16.3090 ;
      RECT 0.0000 10.6960 131.4060 16.3030 ;
      RECT 0.0000 0.0000 19.9780 9.2950 ;
      RECT 0.0000 0.0000 19.9780 9.2950 ;
      RECT 0.0000 0.8000 22.2680 9.2950 ;
      RECT 0.0000 0.8000 22.2680 9.2950 ;
      RECT 0.0000 0.8000 22.2680 0.8020 ;
      RECT 0.8000 10.6950 131.4060 16.3030 ;
      RECT 0.8000 10.6950 131.4060 16.3030 ;
      RECT 0.8000 10.6950 131.4060 16.3030 ;
      RECT 0.8000 10.6950 131.4060 10.6960 ;
      RECT 0.8000 9.2960 130.6060 10.6950 ;
      RECT 0.0000 116.3040 130.6060 116.3130 ;
      RECT 0.0000 41.9680 130.6060 116.3130 ;
      RECT 0.0000 41.9680 130.6060 116.3130 ;
      RECT 0.0000 41.9680 130.6060 116.3130 ;
      RECT 0.0000 41.9680 131.4060 116.3040 ;
      RECT 0.0000 41.9530 130.6060 116.3040 ;
      RECT 0.0000 41.9530 130.6060 116.3040 ;
      RECT 0.0000 41.9530 130.6060 116.3040 ;
      RECT 0.0000 41.9530 130.6060 41.9680 ;
      RECT 0.8000 40.5680 130.6060 41.9530 ;
      RECT 0.0000 18.2430 131.4060 40.5530 ;
      RECT 0.8000 18.2430 130.6060 41.9530 ;
      RECT 0.8000 18.2430 130.6060 41.9530 ;
      RECT 0.8000 18.2430 130.6060 41.9530 ;
      RECT 0.8000 40.5530 131.4060 40.5680 ;
      RECT 0.8000 18.2430 131.4060 40.5680 ;
      RECT 0.8000 18.2430 131.4060 40.5680 ;
      RECT 0.8000 18.2430 131.4060 40.5680 ;
      RECT 0.8000 18.1650 131.4060 40.5530 ;
      RECT 0.8000 18.1650 131.4060 40.5530 ;
      RECT 0.8000 18.1650 131.4060 40.5530 ;
      RECT 0.8000 18.1650 131.4060 18.2430 ;
      RECT 0.8000 16.3090 130.6060 18.1650 ;
      RECT 0.8000 116.3130 130.6060 117.7040 ;
      RECT 0.8000 41.9680 130.6060 117.7040 ;
      RECT 0.8000 41.9680 130.6060 117.7040 ;
      RECT 0.8000 41.9680 130.6060 117.7040 ;
      RECT 0.0000 9.2950 130.6060 9.2960 ;
      RECT 0.0000 0.8020 130.6060 9.2960 ;
      RECT 0.0000 0.8020 130.6060 9.2960 ;
      RECT 0.0000 0.8020 130.6060 9.2960 ;
      RECT 0.0000 0.8020 131.4060 9.2950 ;
    LAYER PO ;
      RECT 0.0000 0.0000 131.4060 154.6780 ;
    LAYER M2 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 40.4530 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 18.3430 ;
      RECT 0.0000 9.1950 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 131.4060 9.1950 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 0.9020 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 135.4590 131.4060 141.1340 ;
      RECT 0.9000 135.4340 131.4060 141.1340 ;
      RECT 0.9000 132.3380 130.5060 141.1340 ;
      RECT 0.9000 135.4340 131.4060 135.4590 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 145.6800 ;
      RECT 0.9000 143.7510 130.5060 144.0800 ;
      RECT 0.0000 148.9090 131.4060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 145.7050 130.5060 148.9090 ;
      RECT 66.8340 0.9000 67.0040 0.9020 ;
      RECT 0.0000 138.1550 130.5060 141.1560 ;
      RECT 0.0000 145.6800 1.5010 147.3090 ;
      RECT 0.0000 142.7560 0.9000 144.0800 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 66.8340 0.9000 67.0040 1.0510 ;
      RECT 128.4050 148.8320 131.4060 148.9090 ;
      RECT 129.9050 145.7050 131.4060 147.2320 ;
      RECT 130.5060 142.7340 131.4060 143.7510 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 132.3080 130.5060 132.3380 ;
      RECT 0.9000 132.3380 130.5060 135.4340 ;
      RECT 0.0000 16.2030 130.5060 16.2090 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 0.9020 ;
      RECT 0.0000 126.6240 130.5060 132.3380 ;
      RECT 0.0000 126.6240 131.4060 132.3080 ;
      RECT 0.9000 126.6240 130.5060 135.4340 ;
      RECT 0.9000 126.6070 131.4060 132.3080 ;
      RECT 0.9000 123.5060 130.5060 132.3080 ;
      RECT 0.9000 126.6070 131.4060 126.6240 ;
      RECT 0.9000 123.5060 130.5060 126.6070 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 10.7960 ;
      RECT 0.9000 9.1960 130.5060 10.7950 ;
      RECT 0.0000 123.4850 130.5060 123.5060 ;
      RECT 0.0000 117.8130 130.5060 123.5060 ;
      RECT 0.0000 117.8130 131.4060 123.4850 ;
      RECT 0.9000 117.8130 130.5060 126.6070 ;
      RECT 0.0000 116.2040 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 131.4060 116.2040 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 117.8130 ;
      RECT 0.9000 116.2130 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 16.2090 130.5060 18.2650 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 42.0680 ;
      RECT 0.0000 18.3430 131.4060 40.4530 ;
      RECT 0.9000 40.4680 130.5060 42.0530 ;
    LAYER M3 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 131.4060 116.2040 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 117.8130 ;
      RECT 0.9000 116.2130 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 16.2090 130.5060 18.2650 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 42.0680 ;
      RECT 0.0000 18.3430 131.4060 40.4530 ;
      RECT 0.9000 40.4680 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 40.4530 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 18.3430 ;
      RECT 0.0000 9.1950 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 131.4060 9.1950 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 0.9020 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 135.4590 131.4060 141.1340 ;
      RECT 0.9000 135.4340 131.4060 141.1340 ;
      RECT 0.9000 132.3380 130.5060 141.1340 ;
      RECT 0.9000 135.4340 131.4060 135.4590 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 145.6800 ;
      RECT 0.9000 143.7510 130.5060 144.0800 ;
      RECT 0.0000 148.9090 131.4060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 145.7050 130.5060 148.9090 ;
      RECT 66.8340 0.9000 67.0040 0.9020 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 138.1550 130.5060 141.1560 ;
      RECT 0.0000 145.6800 1.5010 147.3090 ;
      RECT 0.0000 142.7560 0.9000 144.0800 ;
      RECT 66.8340 0.9000 67.0040 1.0510 ;
      RECT 128.4050 148.8320 131.4060 148.9090 ;
      RECT 129.9050 145.7050 131.4060 147.2320 ;
      RECT 130.5060 142.7340 131.4060 143.7510 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 132.3080 130.5060 132.3380 ;
      RECT 0.9000 132.3380 130.5060 135.4340 ;
      RECT 0.0000 16.2030 130.5060 16.2090 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 0.9020 ;
      RECT 0.0000 126.6240 130.5060 132.3380 ;
      RECT 0.0000 126.6240 131.4060 132.3080 ;
      RECT 0.9000 126.6240 130.5060 135.4340 ;
      RECT 0.9000 126.6070 131.4060 132.3080 ;
      RECT 0.9000 123.5060 130.5060 132.3080 ;
      RECT 0.9000 126.6070 131.4060 126.6240 ;
      RECT 0.9000 123.5060 130.5060 126.6070 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 10.7960 ;
      RECT 0.9000 9.1960 130.5060 10.7950 ;
      RECT 0.0000 123.4850 130.5060 123.5060 ;
      RECT 0.0000 117.8130 130.5060 123.5060 ;
      RECT 0.0000 117.8130 131.4060 123.4850 ;
      RECT 0.9000 117.8130 130.5060 126.6070 ;
      RECT 0.0000 116.2040 130.5060 116.2130 ;
    LAYER M4 ;
      RECT 0.9000 126.6240 130.5060 135.4340 ;
      RECT 0.9000 126.6070 131.4060 132.3080 ;
      RECT 0.9000 123.5060 130.5060 132.3080 ;
      RECT 0.9000 126.6070 131.4060 126.6240 ;
      RECT 0.9000 123.5060 130.5060 126.6070 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 10.7960 ;
      RECT 0.9000 9.1960 130.5060 10.7950 ;
      RECT 0.0000 123.4850 130.5060 123.5060 ;
      RECT 0.0000 117.8130 130.5060 123.5060 ;
      RECT 0.0000 117.8130 131.4060 123.4850 ;
      RECT 0.9000 117.8130 130.5060 126.6070 ;
      RECT 0.0000 116.2040 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 130.5060 116.2130 ;
      RECT 0.0000 42.0680 131.4060 116.2040 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 123.4850 ;
      RECT 0.9000 117.8040 131.4060 117.8130 ;
      RECT 0.9000 116.2130 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 42.0680 130.5060 117.8040 ;
      RECT 0.9000 16.2090 130.5060 18.2650 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 42.0680 ;
      RECT 0.0000 18.3430 131.4060 40.4530 ;
      RECT 0.9000 40.4680 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 40.4530 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 18.3430 ;
      RECT 0.0000 9.1950 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 131.4060 9.1950 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 0.9020 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
      RECT 0.0000 135.4590 131.4060 141.1340 ;
      RECT 0.9000 135.4340 131.4060 141.1340 ;
      RECT 0.9000 132.3380 130.5060 141.1340 ;
      RECT 0.9000 135.4340 131.4060 135.4590 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 147.2320 ;
      RECT 0.9000 141.1560 130.5060 145.6800 ;
      RECT 0.9000 143.7510 130.5060 144.0800 ;
      RECT 0.0000 148.9090 131.4060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 144.0800 130.5060 154.6780 ;
      RECT 0.9000 145.7050 130.5060 148.9090 ;
      RECT 66.8340 0.9000 67.0040 0.9020 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 138.1550 130.5060 141.1560 ;
      RECT 0.0000 145.6800 1.5010 147.3090 ;
      RECT 0.0000 142.7560 0.9000 144.0800 ;
      RECT 66.8340 0.9000 67.0040 1.0510 ;
      RECT 128.4050 148.8320 131.4060 148.9090 ;
      RECT 129.9050 145.7050 131.4060 147.2320 ;
      RECT 130.5060 142.7340 131.4060 143.7510 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 132.3080 130.5060 132.3380 ;
      RECT 0.9000 132.3380 130.5060 135.4340 ;
      RECT 0.0000 16.2030 130.5060 16.2090 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 0.9020 ;
      RECT 0.0000 126.6240 130.5060 132.3380 ;
      RECT 0.0000 126.6240 131.4060 132.3080 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 131.4060 154.6780 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 131.4060 154.6780 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 131.4060 154.6780 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 131.4060 154.6780 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 131.4060 154.6780 ;
    LAYER M5 ;
      RECT 66.8340 0.9000 67.0040 0.9020 ;
      RECT 131.1530 153.6780 131.4060 154.6780 ;
      RECT 0.0000 153.6780 0.3080 154.6780 ;
      RECT 21.4780 0.0000 22.1680 0.9000 ;
      RECT 0.0000 145.7050 1.5010 147.2320 ;
      RECT 0.0000 145.6800 0.9000 145.7050 ;
      RECT 0.0000 147.2320 0.9000 147.3090 ;
      RECT 0.0000 142.7560 0.9000 144.0800 ;
      RECT 0.9000 141.1560 130.5060 142.7340 ;
      RECT 0.9000 142.7340 131.4060 142.7560 ;
      RECT 66.8340 0.9000 67.0040 1.0510 ;
      RECT 129.9050 145.7050 131.4060 147.2320 ;
      RECT 130.5060 142.7560 131.4060 143.7510 ;
      RECT 0.0000 0.0000 19.8780 0.9000 ;
      RECT 0.0000 141.1340 130.5060 141.1560 ;
      RECT 0.0000 42.0680 131.4060 116.2040 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.0000 19.8780 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 9.1950 ;
      RECT 0.0000 0.9000 22.1680 0.9020 ;
      RECT 0.0000 16.2030 130.5060 16.2090 ;
      RECT 0.0000 116.2040 130.5060 116.2130 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 130.5060 16.2090 ;
      RECT 0.0000 10.7960 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 16.2030 ;
      RECT 0.9000 10.7950 131.4060 10.7960 ;
      RECT 0.9000 9.1960 130.5060 10.7950 ;
      RECT 0.9000 143.7510 130.5060 144.0800 ;
      RECT 0.9000 142.7560 130.5060 143.7510 ;
      RECT 0.9000 16.2090 130.5060 18.2650 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 116.2040 ;
      RECT 0.0000 42.0530 130.5060 42.0680 ;
      RECT 0.0000 18.3430 131.4060 40.4530 ;
      RECT 0.9000 40.4680 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 18.3430 130.5060 42.0530 ;
      RECT 0.9000 40.4530 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.3430 131.4060 40.4680 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 40.4530 ;
      RECT 0.9000 18.2650 131.4060 18.3430 ;
      RECT 0.9000 117.8040 131.4060 117.8130 ;
      RECT 0.9000 116.2130 130.5060 117.8040 ;
      RECT 0.0000 148.9090 131.4060 153.6780 ;
      RECT 0.9000 148.8320 131.4060 148.9090 ;
      RECT 0.9000 145.7050 130.5060 148.9090 ;
      RECT 0.9000 147.2320 130.5060 147.3090 ;
      RECT 0.9000 145.7050 130.5060 147.2320 ;
      RECT 0.9000 144.0800 130.5060 147.2320 ;
      RECT 0.9000 144.0800 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 143.7510 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.9000 142.7560 130.5060 147.2320 ;
      RECT 0.0000 135.4590 131.4060 141.1340 ;
      RECT 0.0000 132.3080 130.5060 132.3380 ;
      RECT 0.9000 135.4340 131.4060 135.4590 ;
      RECT 0.9000 132.3380 130.5060 135.4590 ;
      RECT 0.9000 132.3380 130.5060 135.4340 ;
      RECT 0.9000 132.3080 130.5060 135.4340 ;
      RECT 0.0000 126.6240 131.4060 132.3080 ;
      RECT 0.0000 123.4850 130.5060 123.5060 ;
      RECT 0.0000 117.8130 131.4060 123.4850 ;
      RECT 0.9000 126.6070 131.4060 126.6240 ;
      RECT 0.9000 123.5060 130.5060 126.6240 ;
      RECT 0.9000 123.5060 130.5060 126.6070 ;
      RECT 0.9000 123.4850 130.5060 126.6070 ;
      RECT 0.0000 9.1950 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 130.5060 9.1960 ;
      RECT 0.0000 0.9020 131.4060 9.1950 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 0.9000 0.9020 130.5060 16.2030 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 9.1950 ;
      RECT 111.0120 0.9000 131.4060 0.9020 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 9.1950 ;
      RECT 111.5180 0.0000 131.4060 0.9000 ;
  END
END SRAMLP2RW128x32

MACRO SRAMLP1RW32x50
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 90.865 BY 96.244 ;
  SYMMETRY X Y R90 ;

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[18]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[39]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[29]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[37]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[31]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[38]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[16]

  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[46]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[27]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 17.2900 90.8650 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 17.2900 90.8650 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 17.2900 90.8650 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 17.2900 90.8650 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 17.2900 90.8650 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 61.4040 90.8650 61.6040 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 61.4040 90.8650 61.6040 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 61.4040 90.8650 61.6040 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 61.4040 90.8650 61.6040 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 61.4040 90.8650 61.6040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 16.8280 90.8650 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 16.8280 90.8650 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 16.8280 90.8650 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 16.8280 90.8650 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 16.8280 90.8650 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[25]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[12]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[19]

  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[46]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[22]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 70.2240 90.8650 70.4240 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 70.2240 90.8650 70.4240 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 70.2240 90.8650 70.4240 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 70.2240 90.8650 70.4240 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 70.2240 90.8650 70.4240 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 79.0440 90.8650 79.2440 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 79.0440 90.8650 79.2440 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 79.0440 90.8650 79.2440 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 79.0440 90.8650 79.2440 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 79.0440 90.8650 79.2440 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6710 89.4400 90.8650 89.6400 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6710 89.4400 90.8650 89.6400 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6710 89.4400 90.8650 89.6400 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6710 89.4400 90.8650 89.6400 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6710 89.4400 90.8650 89.6400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 62.9940 90.8650 63.1940 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 62.9940 90.8650 63.1940 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 62.9940 90.8650 63.1940 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 62.9940 90.8650 63.1940 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 62.9940 90.8650 63.1940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 71.8140 90.8650 72.0140 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 71.8140 90.8650 72.0140 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 71.8140 90.8650 72.0140 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 71.8140 90.8650 72.0140 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 71.8140 90.8650 72.0140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 89.2000 95.9430 89.4990 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.3010 95.9430 88.6010 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.0010 95.9430 1.3020 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9010 95.9430 2.2020 96.2430 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 77.0510 95.9430 77.3500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.6510 95.9430 44.9500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2520 95.9430 12.5510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.5510 95.9430 72.8500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.1510 95.9430 40.4500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7520 95.9430 8.0510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.3510 95.9430 74.6510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.9510 95.9430 42.2510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5520 95.9430 9.8520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.4520 95.9430 73.7530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.0520 95.9430 41.3530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6530 95.9430 8.9540 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.7520 95.9430 89.0520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.1520 95.9430 85.4520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.3510 95.9430 83.6510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.5510 95.9430 63.8510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.9520 95.9430 60.2520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.3520 95.9430 56.6520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.7520 95.9430 53.0520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.9510 95.9430 51.2510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1520 95.9430 31.4520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5530 95.9430 27.8530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9530 95.9430 24.2530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3530 95.9430 20.6530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5520 95.9430 18.8520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.8510 95.9430 88.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.9510 95.9430 87.2510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.0510 95.9430 86.3510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.2510 95.9430 84.5510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.4500 95.9430 64.7500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.6500 95.9430 62.9500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.7510 95.9430 62.0510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.8510 95.9430 61.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.0510 95.9430 59.3510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.1510 95.9430 58.4510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.2510 95.9430 57.5510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.4510 95.9430 55.7510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.5510 95.9430 54.8510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.6510 95.9430 53.9510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.8510 95.9430 52.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0510 95.9430 32.3510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2510 95.9430 30.5510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3520 95.9430 29.6520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4520 95.9430 28.7520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6520 95.9430 26.9520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7520 95.9430 26.0520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8520 95.9430 25.1520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0520 95.9430 23.3520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1520 95.9430 22.4520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2520 95.9430 21.5520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4520 95.9430 19.7520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1530 95.9430 13.4540 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.8510 95.9430 70.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.5530 95.9430 0.8530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.9520 95.9430 33.2520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.3520 95.9430 65.6520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4530 95.9430 1.7520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.8520 95.9430 34.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.4510 95.9430 37.7510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0520 95.9430 5.3520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.0510 95.9430 68.3520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.6510 95.9430 35.9520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2520 95.9430 3.5530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.9510 95.9430 69.2520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.5510 95.9430 36.8520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.1520 95.9430 4.4530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.7510 95.9430 71.0510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.3510 95.9430 38.6510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9520 95.9430 6.2520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.7510 95.9430 80.0510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.3510 95.9430 47.6510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9520 95.9430 15.2520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.5510 95.9430 81.8500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.1510 95.9430 49.4500 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7520 95.9430 17.0510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.6520 95.9430 80.9520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.2520 95.9430 48.5520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8530 95.9430 16.1530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.1520 95.9430 67.4510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.7520 95.9430 35.0510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3530 95.9430 2.6520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.2510 95.9430 75.5510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.8510 95.9430 43.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4520 95.9430 10.7520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.8510 95.9430 79.1510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.4510 95.9430 46.7510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0520 95.9430 14.3520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.4520 95.9430 82.7530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.0520 95.9430 50.3530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6530 95.9430 17.9540 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.6520 95.9430 71.9520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.2520 95.9430 39.5520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8530 95.9430 7.1530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.1520 95.9430 76.4520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.7520 95.9430 44.0520 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3530 95.9430 11.6530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.9520 95.9430 78.2530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.5520 95.9430 45.8530 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.2520 95.9430 66.5510 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.6510 95.9440 89.9510 96.2440 ;
    END
  END VSS

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6710 86.2410 90.8650 86.4410 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6710 86.2410 90.8650 86.4410 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6710 86.2410 90.8650 86.4410 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6710 86.2410 90.8650 86.4410 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6710 86.2410 90.8650 86.4410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6710 85.8980 90.8650 86.0980 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6710 85.8980 90.8650 86.0980 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6710 85.8980 90.8650 86.0980 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6710 85.8980 90.8650 86.0980 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6710 85.8980 90.8650 86.0980 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.9970 0.0000 70.1970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.9970 0.0000 70.1970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.9970 0.0000 70.1970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.9970 0.0000 70.1970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.9970 0.0000 70.1970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[45]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[3]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[15]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[17]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[32]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[1]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[35]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[23]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.8020 95.9430 3.1020 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.7020 95.9430 4.0020 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.5000 95.9430 86.7990 96.2430 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.4010 95.9430 87.7000 96.2430 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[0]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[9]

  PIN O[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[49]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[34]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[11]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9750 0.0010 3.1750 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9750 0.0010 3.1750 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN I[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[49]

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[44]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[13]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[10]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[10]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[33]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[22]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[8]

  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[47]

  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[47]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[26]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[4]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[42]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[28]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[13]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[36]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[28]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[30]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.694437 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.694437 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9861 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[21]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.648957 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.648957 LAYER M3 ;
    ANTENNAMAXAREACAR 79.77003 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[27]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[24]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[26]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[7]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[40]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[21]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[39]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[14]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[37]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.648957 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.648957 LAYER M3 ;
    ANTENNAMAXAREACAR 79.77003 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[12]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[34]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[1]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[42]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[41]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[30]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[2]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[4]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[43]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[41]

  PIN O[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[48]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[6]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.648957 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.648957 LAYER M3 ;
    ANTENNAMAXAREACAR 79.77003 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[24]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.6650 9.8200 90.8650 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.6650 9.8200 90.8650 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.6650 9.8200 90.8650 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.6650 9.8200 90.8650 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.6650 9.8200 90.8650 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1705 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1705 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.57186 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.57186 LAYER M2 ;
    ANTENNAMAXAREACAR 11.79713 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.52312 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52312 LAYER M3 ;
    ANTENNAMAXAREACAR 15.37747 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.52312 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52312 LAYER M4 ;
    ANTENNAMAXAREACAR 18.95773 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 19.99413 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.694437 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.694437 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9861 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[40]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[20]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.56835 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56835 LAYER M3 ;
  END O[5]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[6]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[19]

  PIN I[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.588357 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.588357 LAYER M3 ;
    ANTENNAMAXAREACAR 76.88431 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[48]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17032 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17032 LAYER M2 ;
    ANTENNAGATEAREA 0.045 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.695457 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.695457 LAYER M3 ;
    ANTENNAMAXAREACAR 106.9737 LAYER M3 ;
    ANTENNAGATEAREA 0.045 LAYER M4 ;
    ANTENNAGATEAREA 0.045 LAYER M5 ;
    ANTENNAGATEAREA 0.045 LAYER M6 ;
    ANTENNAGATEAREA 0.045 LAYER M7 ;
    ANTENNAGATEAREA 0.045 LAYER M8 ;
    ANTENNAGATEAREA 0.045 LAYER M9 ;
    ANTENNAGATEAREA 0.045 LAYER MRDL ;
  END I[2]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.8000 90.0650 96.2440 ;
      RECT 0.0000 0.8000 90.0650 96.2440 ;
      RECT 0.0000 85.2980 90.0710 90.2400 ;
      RECT 0.0000 79.8440 90.8650 85.2980 ;
      RECT 0.0000 78.4440 90.0650 79.8440 ;
      RECT 90.0650 71.0240 90.8650 71.2140 ;
      RECT 90.0650 62.2040 90.8650 62.3940 ;
      RECT 0.0000 0.0000 1.0070 0.8000 ;
      RECT 89.3640 87.0410 90.8650 88.8400 ;
      RECT 0.0000 72.6140 90.8650 78.4440 ;
      RECT 0.0000 69.6240 90.0650 72.6140 ;
      RECT 0.0000 63.7940 90.8650 69.6240 ;
      RECT 0.0000 60.8040 90.0650 63.7940 ;
      RECT 0.0000 18.0900 90.8650 60.8040 ;
      RECT 0.0000 16.2280 90.0650 18.0900 ;
      RECT 0.0000 10.6200 90.8650 16.2280 ;
      RECT 0.0000 9.2200 90.0650 10.6200 ;
      RECT 0.0000 0.8000 90.8650 9.2200 ;
      RECT 70.7970 0.0000 90.8650 9.2200 ;
      RECT 70.7970 0.0000 90.8650 0.8000 ;
      RECT 0.0000 90.2400 90.8650 96.2440 ;
      RECT 0.0000 79.8440 90.0710 96.2440 ;
      RECT 0.0000 0.8000 90.0650 96.2440 ;
      RECT 0.0000 0.8000 90.0650 96.2440 ;
      RECT 0.0000 0.8000 90.0650 96.2440 ;
    LAYER PO ;
      RECT 0.0000 0.0000 90.8650 96.2440 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 90.8650 96.2440 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 90.8650 96.2440 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 90.8650 96.2440 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 90.8650 96.2440 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 90.8650 96.2440 ;
    LAYER M5 ;
      RECT 90.6510 95.2440 90.8650 96.2440 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 90.1990 95.2430 90.8650 95.2440 ;
      RECT 0.0000 0.9000 2.2750 0.9010 ;
      RECT 0.0000 0.9000 2.2750 2.4010 ;
      RECT 89.3640 87.1410 90.8650 88.7400 ;
      RECT 90.1990 94.9430 90.8650 95.2440 ;
      RECT 70.8970 0.0000 90.8650 0.9000 ;
      RECT 0.0000 72.7140 90.8650 78.3440 ;
      RECT 0.0000 69.5240 89.9650 72.7140 ;
      RECT 0.0000 63.8940 90.8650 69.5240 ;
      RECT 0.0000 60.7040 89.9650 63.8940 ;
      RECT 0.0000 18.1900 90.8650 60.7040 ;
      RECT 0.0000 16.1280 89.9650 18.1900 ;
      RECT 0.0000 10.7200 90.8650 16.1280 ;
      RECT 0.0000 9.1200 89.9650 10.7200 ;
      RECT 0.0000 0.9010 90.8650 9.1200 ;
      RECT 3.8750 0.9000 90.8650 9.1200 ;
      RECT 3.8750 0.9000 90.8650 0.9010 ;
      RECT 70.8970 0.0000 90.8650 9.1200 ;
      RECT 0.0000 90.3400 90.8650 95.2430 ;
      RECT 0.0000 79.9440 89.9710 95.2430 ;
      RECT 0.0000 0.9010 89.9650 95.2430 ;
      RECT 0.0000 0.9010 89.9650 95.2430 ;
      RECT 0.0000 0.9010 89.9650 95.2430 ;
      RECT 0.0000 0.9010 89.9650 95.2430 ;
      RECT 0.0000 0.9010 89.9650 95.2430 ;
      RECT 0.0000 85.1980 89.9710 90.3400 ;
      RECT 0.0000 79.9440 90.8650 85.1980 ;
      RECT 0.0000 78.3440 89.9650 79.9440 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 0.0000 0.9000 2.2750 2.4010 ;
      RECT 89.3640 87.1410 90.8650 88.7400 ;
      RECT 70.8970 0.0000 90.8650 0.9000 ;
      RECT 0.0000 72.7140 90.8650 78.3440 ;
      RECT 0.0000 69.5240 89.9650 72.7140 ;
      RECT 0.0000 63.8940 90.8650 69.5240 ;
      RECT 0.0000 60.7040 89.9650 63.8940 ;
      RECT 0.0000 18.1900 90.8650 60.7040 ;
      RECT 0.0000 16.1280 89.9650 18.1900 ;
      RECT 0.0000 10.7200 90.8650 16.1280 ;
      RECT 0.0000 9.1200 89.9650 10.7200 ;
      RECT 0.0000 0.9010 90.8650 9.1200 ;
      RECT 3.8750 0.9000 90.8650 9.1200 ;
      RECT 3.8750 0.9000 90.8650 0.9010 ;
      RECT 70.8970 0.0000 90.8650 9.1200 ;
      RECT 0.0000 90.3400 90.8650 96.2440 ;
      RECT 0.0000 79.9440 89.9710 96.2440 ;
      RECT 0.0000 0.9010 89.9650 96.2440 ;
      RECT 0.0000 0.9010 89.9650 96.2440 ;
      RECT 0.0000 0.9010 89.9650 96.2440 ;
      RECT 0.0000 0.9010 89.9650 96.2440 ;
      RECT 0.0000 0.9010 89.9650 96.2440 ;
      RECT 0.0000 85.1980 89.9710 90.3400 ;
      RECT 0.0000 79.9440 90.8650 85.1980 ;
      RECT 0.0000 78.3440 89.9650 79.9440 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 89.3640 87.1410 90.8650 88.7400 ;
      RECT 0.0000 72.7140 90.8650 78.3440 ;
      RECT 0.0000 69.5240 89.9650 72.7140 ;
      RECT 0.0000 63.8940 90.8650 69.5240 ;
      RECT 0.0000 60.7040 89.9650 63.8940 ;
      RECT 0.0000 18.1900 90.8650 60.7040 ;
      RECT 0.0000 16.1280 89.9650 18.1900 ;
      RECT 0.0000 10.7200 90.8650 16.1280 ;
      RECT 0.0000 9.1200 89.9650 10.7200 ;
      RECT 0.0000 0.9000 90.8650 9.1200 ;
      RECT 70.8970 0.0000 90.8650 9.1200 ;
      RECT 70.8970 0.0000 90.8650 0.9000 ;
      RECT 0.0000 90.3400 90.8650 96.2440 ;
      RECT 0.0000 79.9440 89.9710 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 85.1980 89.9710 90.3400 ;
      RECT 0.0000 79.9440 90.8650 85.1980 ;
      RECT 0.0000 78.3440 89.9650 79.9440 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 89.3640 87.1410 90.8650 88.7400 ;
      RECT 0.0000 72.7140 90.8650 78.3440 ;
      RECT 0.0000 69.5240 89.9650 72.7140 ;
      RECT 0.0000 63.8940 90.8650 69.5240 ;
      RECT 0.0000 60.7040 89.9650 63.8940 ;
      RECT 0.0000 18.1900 90.8650 60.7040 ;
      RECT 0.0000 16.1280 89.9650 18.1900 ;
      RECT 0.0000 10.7200 90.8650 16.1280 ;
      RECT 0.0000 9.1200 89.9650 10.7200 ;
      RECT 0.0000 0.9000 90.8650 9.1200 ;
      RECT 70.8970 0.0000 90.8650 9.1200 ;
      RECT 70.8970 0.0000 90.8650 0.9000 ;
      RECT 0.0000 90.3400 90.8650 96.2440 ;
      RECT 0.0000 79.9440 89.9710 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 0.9000 89.9650 96.2440 ;
      RECT 0.0000 85.1980 89.9710 90.3400 ;
      RECT 0.0000 79.9440 90.8650 85.1980 ;
      RECT 0.0000 78.3440 89.9650 79.9440 ;
  END
END SRAMLP1RW32x50

MACRO SRAMLP1RW64x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 33.296 BY 145.366 ;
  SYMMETRY X Y R90 ;

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.094192 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.094192 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[7]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 16.9030 33.2960 17.1030 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 16.9030 33.2960 17.1030 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 16.9030 33.2960 17.1030 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 16.9030 33.2960 17.1030 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 16.9030 33.2960 17.1030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.093454 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.093454 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[0]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0950 129.1230 33.2950 129.3230 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0950 129.1230 33.2950 129.3230 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0950 129.1230 33.2950 129.3230 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0950 129.1230 33.2950 129.3230 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0950 129.1230 33.2950 129.3230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.094476 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.094476 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[1]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[5]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1010 125.3940 33.2950 125.5940 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1010 125.3940 33.2950 125.5940 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1010 125.3940 33.2950 125.5940 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1010 125.3940 33.2950 125.5940 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1010 125.3940 33.2950 125.5940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 9.8910 33.2960 10.0910 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 9.8910 33.2960 10.0910 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 9.8910 33.2960 10.0910 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 9.8910 33.2960 10.0910 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 9.8910 33.2960 10.0910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 17.3590 33.2960 17.5590 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 17.3590 33.2960 17.5590 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 17.3590 33.2960 17.5590 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 17.3590 33.2960 17.5590 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 17.3590 33.2960 17.5590 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 104.1840 33.2960 104.3840 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 104.1840 33.2960 104.3840 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 104.1840 33.2960 104.3840 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 104.1840 33.2960 104.3840 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 104.1840 33.2960 104.3840 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 111.5460 33.2960 111.7460 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 111.5460 33.2960 111.7460 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 111.5460 33.2960 111.7460 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 111.5460 33.2960 111.7460 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 111.5460 33.2960 111.7460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 113.1040 33.2960 113.3040 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 113.1040 33.2960 113.3040 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 113.1040 33.2960 113.3040 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 113.1040 33.2960 113.3040 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 113.1040 33.2960 113.3040 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 121.8750 33.2960 122.0750 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 121.8750 33.2960 122.0750 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 121.8750 33.2960 122.0750 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 121.8750 33.2960 122.0750 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 121.8750 33.2960 122.0750 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0960 120.3280 33.2960 120.5280 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0960 120.3280 33.2960 120.5280 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0960 120.3280 33.2960 120.5280 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0960 120.3280 33.2960 120.5280 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0960 120.3280 33.2960 120.5280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1010 128.5800 33.2950 128.7800 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1010 128.5800 33.2950 128.7800 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1010 128.5800 33.2950 128.7800 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1010 128.5800 33.2950 128.7800 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1010 128.5800 33.2950 128.7800 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9010 145.0650 29.2000 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.8010 145.0650 30.1000 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.8020 145.0650 3.1020 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.9010 145.0650 2.2020 145.3650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1010 125.0140 33.2950 125.2140 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1010 125.0140 33.2950 125.2140 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1010 125.0140 33.2950 125.2140 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1010 125.0140 33.2950 125.2140 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1010 125.0140 33.2950 125.2140 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    ANTENNADIFFAREA 18.25124 LAYER M1 ;
    ANTENNADIFFAREA 18.25124 LAYER M2 ;
    ANTENNADIFFAREA 18.25124 LAYER M3 ;
    ANTENNADIFFAREA 18.25124 LAYER M4 ;
    ANTENNADIFFAREA 18.25124 LAYER M5 ;
    ANTENNADIFFAREA 18.25124 LAYER M6 ;
    ANTENNADIFFAREA 18.25124 LAYER M7 ;
    ANTENNADIFFAREA 18.25124 LAYER M8 ;
    ANTENNADIFFAREA 18.25124 LAYER M9 ;
    ANTENNADIFFAREA 18.25124 LAYER MRDL ;
    ANTENNAGATEAREA 2.6979 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 32.34852 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 32.34852 LAYER M1 ;
    ANTENNAGATEAREA 2.6979 LAYER M2 ;
    ANTENNAGATEAREA 2.6979 LAYER M3 ;
    ANTENNAGATEAREA 2.6979 LAYER M4 ;
    ANTENNAGATEAREA 2.6979 LAYER M5 ;
    ANTENNAGATEAREA 2.6979 LAYER M6 ;
    ANTENNAGATEAREA 2.6979 LAYER M7 ;
    ANTENNAGATEAREA 2.6979 LAYER M8 ;
    ANTENNAGATEAREA 2.6979 LAYER M9 ;
    ANTENNAGATEAREA 2.6979 LAYER MRDL ;
  END O[3]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 1.0010 145.0650 1.3020 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.1020 145.0650 0.4010 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.6000 145.0660 31.8990 145.3660 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.7010 145.0660 31.0010 145.3660 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.1510 145.0650 4.4520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0510 145.0650 14.3510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4510 145.0650 10.7510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3520 145.0650 2.6510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8520 145.0650 16.1520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7510 145.0650 17.0500 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9510 145.0650 15.2510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6520 145.0650 17.9530 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8520 145.0650 7.1520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3520 145.0650 11.6520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1520 145.0650 13.4530 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2510 145.0650 12.5500 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7510 145.0650 8.0500 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5510 145.0650 9.8510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6520 145.0650 8.9530 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1510 145.0650 31.4510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5520 145.0650 27.8520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9520 145.0650 24.2520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3520 145.0650 20.6520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5510 145.0650 18.8510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0500 145.0650 32.3500 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2500 145.0650 30.5500 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3510 145.0650 29.6510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4510 145.0650 28.7510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6510 145.0650 26.9510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7510 145.0650 26.0510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8510 145.0650 25.1510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0510 145.0650 23.3510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1510 145.0650 22.4510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2510 145.0650 21.5510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4510 145.0650 19.7510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4520 145.0650 1.7510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.5520 145.0650 0.8520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0510 145.0650 5.3510 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2510 145.0650 3.5520 145.3650 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9510 145.0650 6.2510 145.3650 ;
    END
  END VSS

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.094786 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.094786 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[2]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.093762 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.093762 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[4]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.093874 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.093874 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[6]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]
  OBS
    LAYER M1 ;
      RECT 13.3500 0.0000 33.2960 0.8000 ;
      RECT 32.4960 121.1280 33.2960 121.2750 ;
      RECT 32.4960 112.3460 33.2960 112.5040 ;
      RECT 0.0000 0.0000 1.0060 0.8000 ;
      RECT 31.7950 122.6750 33.2960 124.4140 ;
      RECT 31.7950 126.1940 33.2960 127.9800 ;
      RECT 0.0000 129.9230 33.2960 145.3660 ;
      RECT 0.0000 128.5230 32.4950 129.9230 ;
      RECT 0.0000 0.8000 32.4950 129.9230 ;
      RECT 0.0000 122.6750 32.5010 128.5230 ;
      RECT 0.0000 0.8000 32.4960 128.5230 ;
      RECT 0.0000 0.8000 32.4960 128.5230 ;
      RECT 0.0000 0.8000 32.4960 128.5230 ;
      RECT 0.0000 0.8000 32.4960 128.5230 ;
      RECT 0.0000 0.8000 32.4960 128.5230 ;
      RECT 0.0000 119.7280 32.4960 122.6750 ;
      RECT 0.0000 113.9040 33.2960 119.7280 ;
      RECT 0.0000 110.9460 32.4960 113.9040 ;
      RECT 0.0000 104.9840 33.2960 110.9460 ;
      RECT 0.0000 103.5840 32.4960 104.9840 ;
      RECT 0.0000 18.1590 33.2960 103.5840 ;
      RECT 0.0000 16.3030 32.4960 18.1590 ;
      RECT 0.0000 10.6910 33.2960 16.3030 ;
      RECT 0.0000 9.2910 32.4960 10.6910 ;
      RECT 0.0000 0.8000 33.2960 9.2910 ;
      RECT 13.3500 0.0000 33.2960 9.2910 ;
    LAYER PO ;
      RECT 0.0000 0.0000 33.2960 145.3660 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 33.2960 145.3660 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 33.2960 145.3660 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 33.2960 145.3660 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 33.2960 145.3660 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 33.2960 145.3660 ;
    LAYER M5 ;
      RECT 33.0500 144.3650 33.2960 145.3660 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.7950 126.2940 33.2960 127.8800 ;
      RECT 31.7950 122.7750 33.2960 124.3140 ;
      RECT 0.0000 130.0230 33.2960 144.3650 ;
      RECT 0.0000 128.4230 32.3950 130.0230 ;
      RECT 0.0000 0.9000 32.3950 130.0230 ;
      RECT 0.0000 122.7750 32.4010 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 119.6280 32.3960 122.7750 ;
      RECT 0.0000 114.0040 33.2960 119.6280 ;
      RECT 0.0000 110.8460 32.3960 114.0040 ;
      RECT 0.0000 105.0840 33.2960 110.8460 ;
      RECT 0.0000 103.4840 32.3960 105.0840 ;
      RECT 0.0000 18.2590 33.2960 103.4840 ;
      RECT 0.0000 16.2030 32.3960 18.2590 ;
      RECT 0.0000 10.7910 33.2960 16.2030 ;
      RECT 0.0000 9.1910 32.3960 10.7910 ;
      RECT 0.0000 0.9000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 0.9000 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.7950 126.2940 33.2960 127.8800 ;
      RECT 31.7950 122.7750 33.2960 124.3140 ;
      RECT 0.0000 130.0230 33.2960 145.3660 ;
      RECT 0.0000 128.4230 32.3950 130.0230 ;
      RECT 0.0000 0.9000 32.3950 130.0230 ;
      RECT 0.0000 122.7750 32.4010 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 119.6280 32.3960 122.7750 ;
      RECT 0.0000 114.0040 33.2960 119.6280 ;
      RECT 0.0000 110.8460 32.3960 114.0040 ;
      RECT 0.0000 105.0840 33.2960 110.8460 ;
      RECT 0.0000 103.4840 32.3960 105.0840 ;
      RECT 0.0000 18.2590 33.2960 103.4840 ;
      RECT 0.0000 16.2030 32.3960 18.2590 ;
      RECT 0.0000 10.7910 33.2960 16.2030 ;
      RECT 0.0000 9.1910 32.3960 10.7910 ;
      RECT 0.0000 0.9000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 0.9000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.7950 126.2940 33.2960 127.8800 ;
      RECT 31.7950 122.7750 33.2960 124.3140 ;
      RECT 0.0000 130.0230 33.2960 145.3660 ;
      RECT 0.0000 128.4230 32.3950 130.0230 ;
      RECT 0.0000 0.9000 32.3950 130.0230 ;
      RECT 0.0000 122.7750 32.4010 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 119.6280 32.3960 122.7750 ;
      RECT 0.0000 114.0040 33.2960 119.6280 ;
      RECT 0.0000 110.8460 32.3960 114.0040 ;
      RECT 0.0000 105.0840 33.2960 110.8460 ;
      RECT 0.0000 103.4840 32.3960 105.0840 ;
      RECT 0.0000 18.2590 33.2960 103.4840 ;
      RECT 0.0000 16.2030 32.3960 18.2590 ;
      RECT 0.0000 10.7910 33.2960 16.2030 ;
      RECT 0.0000 9.1910 32.3960 10.7910 ;
      RECT 0.0000 0.9000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 0.9000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.7950 122.7750 33.2960 124.3140 ;
      RECT 31.7950 126.2940 33.2960 127.8800 ;
      RECT 0.0000 130.0230 33.2960 145.3660 ;
      RECT 0.0000 128.4230 32.3950 130.0230 ;
      RECT 0.0000 0.9000 32.3950 130.0230 ;
      RECT 0.0000 122.7750 32.4010 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 0.9000 32.3960 128.4230 ;
      RECT 0.0000 119.6280 32.3960 122.7750 ;
      RECT 0.0000 114.0040 33.2960 119.6280 ;
      RECT 0.0000 110.8460 32.3960 114.0040 ;
      RECT 0.0000 105.0840 33.2960 110.8460 ;
      RECT 0.0000 103.4840 32.3960 105.0840 ;
      RECT 0.0000 18.2590 33.2960 103.4840 ;
      RECT 0.0000 16.2030 32.3960 18.2590 ;
      RECT 0.0000 10.7910 33.2960 16.2030 ;
      RECT 0.0000 9.1910 32.3960 10.7910 ;
      RECT 0.0000 0.9000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 9.1910 ;
      RECT 13.4500 0.0000 33.2960 0.9000 ;
  END
END SRAMLP1RW64x8

MACRO SRAMLP1RW64x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 66.611 BY 143.041 ;
  SYMMETRY X Y R90 ;

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.7230 0.0000 1.9230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.7230 0.0000 1.9230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.7230 0.0000 1.9230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.7230 0.0000 1.9230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.7230 0.0000 1.9230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.3770 0.0000 2.5770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.3770 0.0000 2.5770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.3770 0.0000 2.5770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.3770 0.0000 2.5770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.3770 0.0000 2.5770 0.2000 ;
    END
    ANTENNADIFFAREA 3.55776 LAYER M3 ;
    ANTENNADIFFAREA 3.55776 LAYER M4 ;
    ANTENNADIFFAREA 3.55776 LAYER M5 ;
    ANTENNADIFFAREA 3.55776 LAYER M6 ;
    ANTENNADIFFAREA 3.55776 LAYER M7 ;
    ANTENNADIFFAREA 3.55776 LAYER M8 ;
    ANTENNADIFFAREA 3.55776 LAYER M9 ;
    ANTENNADIFFAREA 3.55776 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
    ANTENNAGATEAREA 0.969 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 12.16946 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.16946 LAYER M3 ;
    ANTENNAMAXAREACAR 23.34902 LAYER M3 ;
    ANTENNAGATEAREA 0.969 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 5.0028 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0028 LAYER M4 ;
    ANTENNAMAXAREACAR 28.51182 LAYER M4 ;
    ANTENNAGATEAREA 0.969 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 5.0028 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0028 LAYER M5 ;
    ANTENNAMAXAREACAR 33.67461 LAYER M5 ;
    ANTENNAGATEAREA 0.969 LAYER M6 ;
    ANTENNAGATEAREA 0.969 LAYER M7 ;
    ANTENNAGATEAREA 0.969 LAYER M8 ;
    ANTENNAGATEAREA 0.969 LAYER M9 ;
    ANTENNAGATEAREA 0.969 LAYER MRDL ;
  END O[16]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.0490 0.0000 42.2490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.0490 0.0000 42.2490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.0490 0.0000 42.2490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.0490 0.0000 42.2490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.0490 0.0000 42.2490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[2]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.7630 0.0000 42.9630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.7630 0.0000 42.9630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.7630 0.0000 42.9630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.7630 0.0000 42.9630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.7630 0.0000 42.9630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.4170 0.0000 43.6170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.4170 0.0000 43.6170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.4170 0.0000 43.6170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.4170 0.0000 43.6170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.4170 0.0000 43.6170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[3]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.1310 0.0000 44.3310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.1310 0.0000 44.3310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.1310 0.0000 44.3310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.1310 0.0000 44.3310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.1310 0.0000 44.3310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7850 0.0000 44.9850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7850 0.0000 44.9850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7850 0.0000 44.9850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7850 0.0000 44.9850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7850 0.0000 44.9850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[5]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4110 9.8910 66.6110 10.0910 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4110 9.8910 66.6110 10.0910 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4110 9.8910 66.6110 10.0910 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4110 9.8910 66.6110 10.0910 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4110 9.8910 66.6110 10.0910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4110 16.9010 66.6110 17.1010 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4110 16.9010 66.6110 17.1010 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4110 16.9010 66.6110 17.1010 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4110 16.9010 66.6110 17.1010 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4110 16.9010 66.6110 17.1010 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4110 17.3630 66.6110 17.5630 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4110 17.3630 66.6110 17.5630 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4110 17.3630 66.6110 17.5630 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4110 17.3630 66.6110 17.5630 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4110 17.3630 66.6110 17.5630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4140 97.8550 66.6110 98.0550 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4140 97.8550 66.6110 98.0550 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4140 97.8550 66.6110 98.0550 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4140 97.8550 66.6110 98.0550 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4140 97.8550 66.6110 98.0550 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4140 105.5720 66.6110 105.7720 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4140 105.5720 66.6110 105.7720 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4140 105.5720 66.6110 105.7720 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4140 105.5720 66.6110 105.7720 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4140 105.5720 66.6110 105.7720 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4120 107.1630 66.6110 107.3630 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4120 107.1630 66.6110 107.3630 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4120 107.1630 66.6110 107.3630 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4120 107.1630 66.6110 107.3630 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4120 107.1630 66.6110 107.3630 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4270 114.3920 66.6110 114.5920 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4270 114.3920 66.6110 114.5920 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4270 114.3920 66.6110 114.5920 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4270 114.3920 66.6110 114.5920 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4270 114.3920 66.6110 114.5920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4140 115.9820 66.6110 116.1820 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4140 115.9820 66.6110 116.1820 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4140 115.9820 66.6110 116.1820 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4140 115.9820 66.6110 116.1820 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4140 115.9820 66.6110 116.1820 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4110 117.4280 66.6110 117.6280 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4110 117.4280 66.6110 117.6280 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4110 117.4280 66.6110 117.6280 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4110 117.4280 66.6110 117.6280 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4110 117.4280 66.6110 117.6280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4170 119.0760 66.6110 119.2760 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4170 119.0760 66.6110 119.2760 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4170 119.0760 66.6110 119.2760 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4170 119.0760 66.6110 119.2760 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4170 119.0760 66.6110 119.2760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4170 119.7400 66.6110 119.9400 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4170 119.7400 66.6110 119.9400 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4170 119.7400 66.6110 119.9400 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4170 119.7400 66.6110 119.9400 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4170 119.7400 66.6110 119.9400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.4170 122.5890 66.6110 122.7890 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.4170 122.5890 66.6110 122.7890 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.4170 122.5890 66.6110 122.7890 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.4170 122.5890 66.6110 122.7890 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.4170 122.5890 66.6110 122.7890 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.4900 0.0000 45.6900 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.4900 0.0000 45.6900 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.4900 0.0000 45.6900 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.4900 0.0000 45.6900 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.4900 0.0000 45.6900 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.3690 0.0000 28.5690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.3690 0.0000 28.5690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.3690 0.0000 28.5690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.3690 0.0000 28.5690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.3690 0.0000 28.5690 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[13]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.0830 0.0000 29.2830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.0830 0.0000 29.2830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.0830 0.0000 29.2830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.0830 0.0000 29.2830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.0830 0.0000 29.2830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.7370 0.0000 29.9370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.7370 0.0000 29.9370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.7370 0.0000 29.9370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.7370 0.0000 29.9370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.7370 0.0000 29.9370 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[6]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.4510 0.0000 30.6510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.4510 0.0000 30.6510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.4510 0.0000 30.6510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.4510 0.0000 30.6510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.4510 0.0000 30.6510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.1050 0.0000 31.3050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.1050 0.0000 31.3050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.1050 0.0000 31.3050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.1050 0.0000 31.3050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.1050 0.0000 31.3050 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[0]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1870 0.0000 33.3870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1870 0.0000 33.3870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1870 0.0000 33.3870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1870 0.0000 33.3870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1870 0.0000 33.3870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.8410 0.0000 34.0410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.8410 0.0000 34.0410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.8410 0.0000 34.0410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.8410 0.0000 34.0410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.8410 0.0000 34.0410 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[8]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.5550 0.0000 34.7550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.5550 0.0000 34.7550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.5550 0.0000 34.7550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.5550 0.0000 34.7550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.5550 0.0000 34.7550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.2090 0.0000 35.4090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.2090 0.0000 35.4090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.2090 0.0000 35.4090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.2090 0.0000 35.4090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.2090 0.0000 35.4090 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[14]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.9230 0.0000 36.1230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.9230 0.0000 36.1230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.9230 0.0000 36.1230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.9230 0.0000 36.1230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.9230 0.0000 36.1230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.5770 0.0000 36.7770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.5770 0.0000 36.7770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.5770 0.0000 36.7770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.5770 0.0000 36.7770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.5770 0.0000 36.7770 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[9]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.2910 0.0000 37.4910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.2910 0.0000 37.4910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.2910 0.0000 37.4910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.2910 0.0000 37.4910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.2910 0.0000 37.4910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.9450 0.0000 38.1450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.9450 0.0000 38.1450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.9450 0.0000 38.1450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.9450 0.0000 38.1450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.9450 0.0000 38.1450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[15]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.6590 0.0000 38.8590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.6590 0.0000 38.8590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.6590 0.0000 38.8590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.6590 0.0000 38.8590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.6590 0.0000 38.8590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.3130 0.0000 39.5130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.3130 0.0000 39.5130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.3130 0.0000 39.5130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.3130 0.0000 39.5130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.3130 0.0000 39.5130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[11]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.0270 0.0000 40.2270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.0270 0.0000 40.2270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.0270 0.0000 40.2270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.0270 0.0000 40.2270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.0270 0.0000 40.2270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.6810 0.0000 40.8810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.6810 0.0000 40.8810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.6810 0.0000 40.8810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.6810 0.0000 40.8810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.6810 0.0000 40.8810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[12]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.3950 0.0000 41.5950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.3950 0.0000 41.5950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.3950 0.0000 41.5950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.3950 0.0000 41.5950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.3950 0.0000 41.5950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.4030 0.0000 15.6030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.4030 0.0000 15.6030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.4030 0.0000 15.6030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.4030 0.0000 15.6030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.4030 0.0000 15.6030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.0570 0.0000 16.2570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.0570 0.0000 16.2570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.0570 0.0000 16.2570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.0570 0.0000 16.2570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.0570 0.0000 16.2570 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[25]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.7710 0.0000 16.9710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.7710 0.0000 16.9710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.7710 0.0000 16.9710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.7710 0.0000 16.9710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.7710 0.0000 16.9710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 17.4250 0.0000 17.6250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.4250 0.0000 17.6250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.4250 0.0000 17.6250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 17.4250 0.0000 17.6250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 17.4250 0.0000 17.6250 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[26]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.1390 0.0000 18.3390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.1390 0.0000 18.3390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.1390 0.0000 18.3390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.1390 0.0000 18.3390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.1390 0.0000 18.3390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.7930 0.0000 18.9930 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.7930 0.0000 18.9930 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.7930 0.0000 18.9930 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.7930 0.0000 18.9930 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.7930 0.0000 18.9930 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[27]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 19.5070 0.0000 19.7070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.5070 0.0000 19.7070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.5070 0.0000 19.7070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.5070 0.0000 19.7070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 19.5070 0.0000 19.7070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.1610 0.0000 20.3610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.1610 0.0000 20.3610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.1610 0.0000 20.3610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.1610 0.0000 20.3610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.1610 0.0000 20.3610 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[28]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.8750 0.0000 21.0750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.8750 0.0000 21.0750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.8750 0.0000 21.0750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.8750 0.0000 21.0750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.8750 0.0000 21.0750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.5290 0.0000 21.7290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.5290 0.0000 21.7290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.5290 0.0000 21.7290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.5290 0.0000 21.7290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.5290 0.0000 21.7290 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[29]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.2430 0.0000 22.4430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.2430 0.0000 22.4430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.2430 0.0000 22.4430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.2430 0.0000 22.4430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.2430 0.0000 22.4430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8970 0.0000 23.0970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8970 0.0000 23.0970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8970 0.0000 23.0970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8970 0.0000 23.0970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8970 0.0000 23.0970 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[30]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.6110 0.0000 23.8110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.6110 0.0000 23.8110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.6110 0.0000 23.8110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.6110 0.0000 23.8110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.6110 0.0000 23.8110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.2650 0.0000 24.4650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.2650 0.0000 24.4650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.2650 0.0000 24.4650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.2650 0.0000 24.4650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.2650 0.0000 24.4650 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[31]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.9790 0.0000 25.1790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.9790 0.0000 25.1790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.9790 0.0000 25.1790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.9790 0.0000 25.1790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.9790 0.0000 25.1790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.6330 0.0000 25.8330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.6330 0.0000 25.8330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.6330 0.0000 25.8330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.6330 0.0000 25.8330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.6330 0.0000 25.8330 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[7]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.3470 0.0000 26.5470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.3470 0.0000 26.5470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.3470 0.0000 26.5470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.3470 0.0000 26.5470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.3470 0.0000 26.5470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.0010 0.0000 27.2010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.0010 0.0000 27.2010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.0010 0.0000 27.2010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.0010 0.0000 27.2010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.0010 0.0000 27.2010 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[4]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.7150 0.0000 27.9150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.7150 0.0000 27.9150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.7150 0.0000 27.9150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.7150 0.0000 27.9150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.7150 0.0000 27.9150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.0910 0.0000 3.2910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.0910 0.0000 3.2910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.0910 0.0000 3.2910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.0910 0.0000 3.2910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.0910 0.0000 3.2910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.7450 0.0000 3.9450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.7450 0.0000 3.9450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.7450 0.0000 3.9450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.7450 0.0000 3.9450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.7450 0.0000 3.9450 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[17]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.4590 0.0000 4.6590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.4590 0.0000 4.6590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.4590 0.0000 4.6590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.4590 0.0000 4.6590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.4590 0.0000 4.6590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.1130 0.0000 5.3130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.1130 0.0000 5.3130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.1130 0.0000 5.3130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.1130 0.0000 5.3130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.1130 0.0000 5.3130 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[18]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.8270 0.0000 6.0270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.8270 0.0000 6.0270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.8270 0.0000 6.0270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.8270 0.0000 6.0270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.8270 0.0000 6.0270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.4810 0.0000 6.6810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.4810 0.0000 6.6810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.4810 0.0000 6.6810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.4810 0.0000 6.6810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.4810 0.0000 6.6810 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[19]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.1950 0.0000 7.3950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.1950 0.0000 7.3950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.1950 0.0000 7.3950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.1950 0.0000 7.3950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.1950 0.0000 7.3950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.8490 0.0000 8.0490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.8490 0.0000 8.0490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.8490 0.0000 8.0490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.8490 0.0000 8.0490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.8490 0.0000 8.0490 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[20]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.5630 0.0000 8.7630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.5630 0.0000 8.7630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.5630 0.0000 8.7630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.5630 0.0000 8.7630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.5630 0.0000 8.7630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.2170 0.0000 9.4170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.2170 0.0000 9.4170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.2170 0.0000 9.4170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.2170 0.0000 9.4170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.2170 0.0000 9.4170 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[21]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.9310 0.0000 10.1310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.9310 0.0000 10.1310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.9310 0.0000 10.1310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.9310 0.0000 10.1310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.9310 0.0000 10.1310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.5850 0.0000 10.7850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.5850 0.0000 10.7850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.5850 0.0000 10.7850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.5850 0.0000 10.7850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.5850 0.0000 10.7850 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[10]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.2990 0.0000 11.4990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.2990 0.0000 11.4990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.2990 0.0000 11.4990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.2990 0.0000 11.4990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.2990 0.0000 11.4990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.9530 0.0000 12.1530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.9530 0.0000 12.1530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.9530 0.0000 12.1530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.9530 0.0000 12.1530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.9530 0.0000 12.1530 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[22]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.6670 0.0000 12.8670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.6670 0.0000 12.8670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.6670 0.0000 12.8670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.6670 0.0000 12.8670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.6670 0.0000 12.8670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.3210 0.0000 13.5210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.3210 0.0000 13.5210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.3210 0.0000 13.5210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.3210 0.0000 13.5210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.3210 0.0000 13.5210 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[23]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.0350 0.0000 14.2350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.0350 0.0000 14.2350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.0350 0.0000 14.2350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.0350 0.0000 14.2350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.0350 0.0000 14.2350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.6890 0.0000 14.8890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.6890 0.0000 14.8890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.6890 0.0000 14.8890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.6890 0.0000 14.8890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.6890 0.0000 14.8890 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[24]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.8190 0.0000 32.0190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.8190 0.0000 32.0190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.8190 0.0000 32.0190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.8190 0.0000 32.0190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.8190 0.0000 32.0190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.3700 142.7410 57.6690 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.2710 142.7410 58.5720 143.0410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.0210 142.7410 56.3220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.8210 142.7410 40.1220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.6210 142.7410 23.9220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.4210 142.7410 7.7220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.6200 142.7410 50.9210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.4200 142.7410 34.7210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.2200 142.7410 18.5210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.0200 142.7410 2.3210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.5200 142.7410 51.8210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.3200 142.7410 35.6210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.1200 142.7410 19.4210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.9200 142.7410 3.2210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.1200 142.7410 55.4190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.9200 142.7410 39.2190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.7200 142.7410 23.0190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.5200 142.7410 6.8190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.4200 142.7410 52.7200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.2200 142.7410 36.5200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.0200 142.7410 20.3200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.8200 142.7410 4.1200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.2210 142.7410 54.5210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.0210 142.7410 38.3210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.8210 142.7410 22.1210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.6210 142.7410 5.9210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.3200 142.7410 53.6200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.1200 142.7410 37.4200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.9200 142.7410 21.2200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.7200 142.7410 5.0200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.7210 142.7410 50.0200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.5210 142.7410 33.8200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.3210 142.7410 17.6200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.1210 142.7410 1.4200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.5210 142.7410 60.8220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.3210 142.7410 44.6220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.1210 142.7410 28.4220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.9210 142.7410 12.2220 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.9200 142.7410 57.2200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.7200 142.7410 41.0200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.5200 142.7410 24.8200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.3200 142.7410 8.6200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.0210 142.7410 65.3200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.8210 142.7410 49.1200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.6210 142.7410 32.9200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.4210 142.7410 16.7200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.2210 142.7410 0.5200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.4200 142.7410 61.7200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.2200 142.7410 45.5200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.0200 142.7410 29.3200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.8200 142.7410 13.1200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.3200 142.7410 62.6200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.1200 142.7410 46.4200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.9200 142.7410 30.2200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.7200 142.7410 14.0200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.7210 142.7410 59.0210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.5210 142.7410 42.8210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.3210 142.7410 26.6210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.1210 142.7410 10.4210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.1210 142.7410 64.4210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.9210 142.7410 48.2210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.7210 142.7410 32.0210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.5210 142.7410 15.8210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.6200 142.7410 59.9190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.4200 142.7410 43.7190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.2200 142.7410 27.5190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.0200 142.7410 11.3190 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.8200 142.7410 58.1200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.6210 142.7410 14.9210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.8210 142.7410 31.1210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.0210 142.7410 47.3210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.2210 142.7410 63.5210 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.2200 142.7410 9.5200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.4200 142.7410 25.7200 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.6200 142.7410 41.9200 143.0410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VSS

  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.6700 142.7410 63.9700 143.0410 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.5700 142.7410 64.8710 143.0410 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDD

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.4730 0.0000 32.6730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.4730 0.0000 32.6730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.4730 0.0000 32.6730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.4730 0.0000 32.6730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.4730 0.0000 32.6730 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.17752 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.17752 LAYER M2 ;
  END O[1]
  OBS
    LAYER M1 ;
      RECT 0.0000 107.9630 65.8270 115.3820 ;
      RECT 0.0000 107.9630 66.6110 113.7920 ;
      RECT 0.0000 106.5630 65.8120 107.9630 ;
      RECT 0.0000 104.9720 65.8140 106.5630 ;
      RECT 0.0000 18.1630 65.8140 106.5630 ;
      RECT 0.0000 18.1630 65.8140 106.5630 ;
      RECT 0.0000 98.6550 66.6110 104.9720 ;
      RECT 0.0000 97.2550 65.8140 98.6550 ;
      RECT 0.0000 18.1630 66.6110 97.2550 ;
      RECT 0.0000 16.3010 65.8110 18.1630 ;
      RECT 0.0000 10.6910 66.6110 16.3010 ;
      RECT 0.0000 9.2910 65.8110 10.6910 ;
      RECT 0.0000 0.8000 66.6110 9.2910 ;
      RECT 46.2900 0.0000 66.6110 9.2910 ;
      RECT 46.2900 0.0000 66.6110 0.8000 ;
      RECT 0.0000 123.3890 66.6110 143.0410 ;
      RECT 0.0000 118.2280 65.8170 143.0410 ;
      RECT 0.0000 0.8000 65.8110 143.0410 ;
      RECT 0.0000 0.8000 65.8110 143.0410 ;
      RECT 0.0000 0.8000 65.8110 143.0410 ;
      RECT 0.0000 118.2280 65.8170 123.3890 ;
      RECT 0.0000 116.8280 65.8110 118.2280 ;
      RECT 65.8140 106.3720 66.6110 106.5630 ;
      RECT 65.8270 115.1920 66.6110 115.3820 ;
      RECT 65.8170 118.2280 66.6110 118.4760 ;
      RECT 0.0000 0.0000 1.1230 0.8000 ;
      RECT 65.8170 120.5400 66.6110 121.9890 ;
      RECT 0.0000 115.3820 65.8140 116.8280 ;
      RECT 0.0000 107.9630 65.8140 116.8280 ;
      RECT 0.0000 18.1630 65.8120 116.8280 ;
      RECT 0.0000 113.7920 65.8270 115.3820 ;
    LAYER PO ;
      RECT 0.0000 0.0000 66.6110 143.0410 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 66.6110 143.0410 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 66.6110 143.0410 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 66.6110 143.0410 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 66.6110 143.0410 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 66.6110 143.0410 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 1.0230 0.9000 ;
      RECT 66.0200 142.0410 66.6110 143.0410 ;
      RECT 65.7170 120.6400 66.6110 121.8890 ;
      RECT 0.0000 115.2820 65.7140 116.7280 ;
      RECT 0.0000 108.0630 65.7140 116.7280 ;
      RECT 0.0000 18.2630 65.7120 116.7280 ;
      RECT 0.0000 113.6920 65.7270 115.2820 ;
      RECT 0.0000 108.0630 65.7270 115.2820 ;
      RECT 0.0000 108.0630 66.6110 113.6920 ;
      RECT 0.0000 106.4630 65.7120 108.0630 ;
      RECT 0.0000 104.8720 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 98.7550 66.6110 104.8720 ;
      RECT 0.0000 97.1550 65.7140 98.7550 ;
      RECT 0.0000 18.2630 66.6110 97.1550 ;
      RECT 0.0000 16.2010 65.7110 18.2630 ;
      RECT 0.0000 10.7910 66.6110 16.2010 ;
      RECT 0.0000 9.1910 65.7110 10.7910 ;
      RECT 0.0000 0.9000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 0.9000 ;
      RECT 0.0000 123.4890 66.6110 142.0410 ;
      RECT 0.0000 118.3280 65.7170 142.0410 ;
      RECT 0.0000 0.9000 65.7110 142.0410 ;
      RECT 0.0000 0.9000 65.7110 142.0410 ;
      RECT 0.0000 0.9000 65.7110 142.0410 ;
      RECT 0.0000 118.3280 65.7170 123.4890 ;
      RECT 0.0000 116.7280 65.7110 118.3280 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1.0230 0.9000 ;
      RECT 65.7170 120.6400 66.6110 121.8890 ;
      RECT 0.0000 115.2820 65.7140 116.7280 ;
      RECT 0.0000 108.0630 65.7140 116.7280 ;
      RECT 0.0000 18.2630 65.7120 116.7280 ;
      RECT 0.0000 113.6920 65.7270 115.2820 ;
      RECT 0.0000 108.0630 65.7270 115.2820 ;
      RECT 0.0000 108.0630 66.6110 113.6920 ;
      RECT 0.0000 106.4630 65.7120 108.0630 ;
      RECT 0.0000 104.8720 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 98.7550 66.6110 104.8720 ;
      RECT 0.0000 97.1550 65.7140 98.7550 ;
      RECT 0.0000 18.2630 66.6110 97.1550 ;
      RECT 0.0000 16.2010 65.7110 18.2630 ;
      RECT 0.0000 10.7910 66.6110 16.2010 ;
      RECT 0.0000 9.1910 65.7110 10.7910 ;
      RECT 0.0000 0.9000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 0.9000 ;
      RECT 0.0000 123.4890 66.6110 143.0410 ;
      RECT 0.0000 118.3280 65.7170 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 118.3280 65.7170 123.4890 ;
      RECT 0.0000 116.7280 65.7110 118.3280 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1.0230 0.9000 ;
      RECT 65.7170 120.6400 66.6110 121.8890 ;
      RECT 0.0000 115.2820 65.7140 116.7280 ;
      RECT 0.0000 108.0630 65.7140 116.7280 ;
      RECT 0.0000 18.2630 65.7120 116.7280 ;
      RECT 0.0000 113.6920 65.7270 115.2820 ;
      RECT 0.0000 108.0630 65.7270 115.2820 ;
      RECT 0.0000 108.0630 66.6110 113.6920 ;
      RECT 0.0000 106.4630 65.7120 108.0630 ;
      RECT 0.0000 104.8720 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 98.7550 66.6110 104.8720 ;
      RECT 0.0000 97.1550 65.7140 98.7550 ;
      RECT 0.0000 18.2630 66.6110 97.1550 ;
      RECT 0.0000 16.2010 65.7110 18.2630 ;
      RECT 0.0000 10.7910 66.6110 16.2010 ;
      RECT 0.0000 9.1910 65.7110 10.7910 ;
      RECT 0.0000 0.9000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 0.9000 ;
      RECT 0.0000 123.4890 66.6110 143.0410 ;
      RECT 0.0000 118.3280 65.7170 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 118.3280 65.7170 123.4890 ;
      RECT 0.0000 116.7280 65.7110 118.3280 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1.0230 0.9000 ;
      RECT 65.7170 120.6400 66.6110 121.8890 ;
      RECT 0.0000 115.2820 65.7140 116.7280 ;
      RECT 0.0000 108.0630 65.7140 116.7280 ;
      RECT 0.0000 18.2630 65.7120 116.7280 ;
      RECT 0.0000 113.6920 65.7270 115.2820 ;
      RECT 0.0000 108.0630 65.7270 115.2820 ;
      RECT 0.0000 108.0630 66.6110 113.6920 ;
      RECT 0.0000 106.4630 65.7120 108.0630 ;
      RECT 0.0000 104.8720 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 18.2630 65.7140 106.4630 ;
      RECT 0.0000 98.7550 66.6110 104.8720 ;
      RECT 0.0000 97.1550 65.7140 98.7550 ;
      RECT 0.0000 18.2630 66.6110 97.1550 ;
      RECT 0.0000 16.2010 65.7110 18.2630 ;
      RECT 0.0000 10.7910 66.6110 16.2010 ;
      RECT 0.0000 9.1910 65.7110 10.7910 ;
      RECT 0.0000 0.9000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 9.1910 ;
      RECT 46.3900 0.0000 66.6110 0.9000 ;
      RECT 0.0000 123.4890 66.6110 143.0410 ;
      RECT 0.0000 118.3280 65.7170 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 0.9000 65.7110 143.0410 ;
      RECT 0.0000 118.3280 65.7170 123.4890 ;
      RECT 0.0000 116.7280 65.7110 118.3280 ;
  END
END SRAMLP1RW64x32

MACRO SRAMLP1RW64x34
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 69.062 BY 142.71 ;
  SYMMETRY X Y R90 ;

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1160 0.0000 9.3160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1160 0.0000 9.3160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1160 0.0000 9.3160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1160 0.0000 9.3160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1160 0.0000 9.3160 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[11]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0120 0.0000 5.2120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0120 0.0000 5.2120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0120 0.0000 5.2120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0120 0.0000 5.2120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0120 0.0000 5.2120 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[32]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8530 0.0000 12.0530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8530 0.0000 12.0530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8530 0.0000 12.0530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8530 0.0000 12.0530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8530 0.0000 12.0530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[13]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.4880 0.0000 10.6880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.4880 0.0000 10.6880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.4880 0.0000 10.6880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.4880 0.0000 10.6880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.4880 0.0000 10.6880 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[12]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 65.0980 142.4100 65.3980 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.1980 142.4100 64.4970 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.1980 142.4100 1.4980 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.2980 142.4100 0.5990 142.7100 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 58.3480 142.4100 58.6480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.5480 142.4100 56.8480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.6480 142.4100 55.9480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.7480 142.4100 55.0480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.9480 142.4100 53.2480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.0480 142.4100 52.3480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.1480 142.4100 51.4480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.3480 142.4100 49.6480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.5480 142.4100 65.8480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.0480 142.4100 61.3480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.4490 142.4100 57.7490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.8490 142.4100 54.1490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.2490 142.4100 50.5490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.4480 142.4100 48.7480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.2480 142.4100 23.5480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.8490 142.4100 27.1480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.0480 142.4100 25.3480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.8480 142.4100 45.1480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.1480 142.4100 42.4470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.9480 142.4100 44.2480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.6480 142.4100 46.9470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.7490 142.4100 46.0490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.0490 142.4100 43.3500 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.5490 142.4100 47.8500 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.9480 142.4100 35.2480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.3490 142.4100 31.6480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.4490 142.4100 30.7490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.4480 142.4100 39.7480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.6480 142.4100 37.9470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.8480 142.4100 36.1480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.7490 142.4100 28.0480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.4490 142.4100 21.7480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.9490 142.4100 26.2490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.7490 142.4100 37.0490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.2490 142.4100 41.5490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.3480 142.4100 40.6480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.2490 142.4100 32.5480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.5490 142.4100 38.8500 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.5480 142.4100 29.8490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.6480 142.4100 28.9490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.5490 142.4100 20.8490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.0480 142.4100 34.3490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.1480 142.4100 33.4490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.1490 142.4100 24.4490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.1480 142.4100 6.4490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.0480 142.4100 7.3490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.6480 142.4100 1.9490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.5480 142.4100 2.8490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.9490 142.4100 8.2490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.2490 142.4100 5.5480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.4490 142.4100 3.7490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.3490 142.4100 4.6480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.7480 142.4100 1.0480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.2480 142.4100 14.5490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.1480 142.4100 15.4490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.0480 142.4100 16.3490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.7480 142.4100 19.0480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.8490 142.4100 18.1490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.9490 142.4100 17.2490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.5480 142.4100 11.8480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.6490 142.4100 10.9490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.8490 142.4100 9.1480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.7480 142.4100 10.0480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.4490 142.4100 12.7480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.3480 142.4100 13.6480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.3480 142.4100 22.6490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.6480 142.4100 19.9490 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.3470 142.4100 67.6470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.2480 142.4100 59.5480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.1470 142.4100 60.4470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.9470 142.4100 62.2470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.8470 142.4100 63.1470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.7480 142.4100 64.0480 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.6470 142.4100 64.9470 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.4470 142.4100 66.7470 142.7100 ;
    END
  END VSS

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 105.2060 69.0620 105.4060 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 105.2060 69.0620 105.4060 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 105.2060 69.0620 105.4060 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 105.2060 69.0620 105.4060 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 105.2060 69.0620 105.4060 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2330 0.0000 26.4330 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2330 0.0000 26.4330 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2330 0.0000 26.4330 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2330 0.0000 26.4330 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2330 0.0000 26.4330 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 16.9940 69.0620 17.1940 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 16.9940 69.0620 17.1940 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 16.9940 69.0620 17.1940 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 16.9940 69.0620 17.1940 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 16.9940 69.0620 17.1940 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 86.5860 69.0620 86.7860 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 86.5860 69.0620 86.7860 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 86.5860 69.0620 86.7860 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 86.5860 69.0620 86.7860 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 86.5860 69.0620 86.7860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1100 0.0000 48.3100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1100 0.0000 48.3100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1100 0.0000 48.3100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1100 0.0000 48.3100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1100 0.0000 48.3100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.1290 0.0000 22.3290 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.1290 0.0000 22.3290 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.1290 0.0000 22.3290 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.1290 0.0000 22.3290 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.1290 0.0000 22.3290 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3800 0.0000 6.5800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3800 0.0000 6.5800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3800 0.0000 6.5800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3800 0.0000 6.5800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3800 0.0000 6.5800 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[33]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8650 0.0000 25.0650 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8650 0.0000 25.0650 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8650 0.0000 25.0650 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8650 0.0000 25.0650 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8650 0.0000 25.0650 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.6010 0.0000 27.8010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.6010 0.0000 27.8010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.6010 0.0000 27.8010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.6010 0.0000 27.8010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.6010 0.0000 27.8010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.7610 0.0000 20.9610 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.7610 0.0000 20.9610 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.7610 0.0000 20.9610 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.7610 0.0000 20.9610 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.7610 0.0000 20.9610 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9690 0.0000 29.1690 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9690 0.0000 29.1690 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9690 0.0000 29.1690 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9690 0.0000 29.1690 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9690 0.0000 29.1690 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3370 0.0000 30.5370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3370 0.0000 30.5370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3370 0.0000 30.5370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3370 0.0000 30.5370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3370 0.0000 30.5370 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7050 0.0000 31.9050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7050 0.0000 31.9050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7050 0.0000 31.9050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7050 0.0000 31.9050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7050 0.0000 31.9050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0730 0.0000 33.2730 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0730 0.0000 33.2730 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0730 0.0000 33.2730 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0730 0.0000 33.2730 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0730 0.0000 33.2730 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4410 0.0000 34.6410 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4410 0.0000 34.6410 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4410 0.0000 34.6410 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4410 0.0000 34.6410 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4410 0.0000 34.6410 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1770 0.0000 37.3770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1770 0.0000 37.3770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1770 0.0000 37.3770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1770 0.0000 37.3770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1770 0.0000 37.3770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8090 0.0000 36.0090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8090 0.0000 36.0090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8090 0.0000 36.0090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8090 0.0000 36.0090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8090 0.0000 36.0090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5450 0.0000 38.7450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5450 0.0000 38.7450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5450 0.0000 38.7450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5450 0.0000 38.7450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5450 0.0000 38.7450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9130 0.0000 40.1130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9130 0.0000 40.1130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9130 0.0000 40.1130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9130 0.0000 40.1130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9130 0.0000 40.1130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2810 0.0000 41.4810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2810 0.0000 41.4810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2810 0.0000 41.4810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2810 0.0000 41.4810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2810 0.0000 41.4810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6490 0.0000 42.8490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6490 0.0000 42.8490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6490 0.0000 42.8490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6490 0.0000 42.8490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6490 0.0000 42.8490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0170 0.0000 44.2170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0170 0.0000 44.2170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0170 0.0000 44.2170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0170 0.0000 44.2170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0170 0.0000 44.2170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3850 0.0030 45.5850 0.2030 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3850 0.0030 45.5850 0.2030 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3850 0.0030 45.5850 0.2030 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3850 0.0030 45.5850 0.2030 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3850 0.0030 45.5850 0.2030 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7530 0.0000 46.9530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7530 0.0000 46.9530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7530 0.0000 46.9530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7530 0.0000 46.9530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7530 0.0000 46.9530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 106.7960 69.0620 106.9960 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 106.7960 69.0620 106.9960 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 106.7960 69.0620 106.9960 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 106.7960 69.0620 106.9960 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 106.7960 69.0620 106.9960 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 97.9760 69.0620 98.1760 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 97.9760 69.0620 98.1760 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 97.9760 69.0620 98.1760 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 97.9760 69.0620 98.1760 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 97.9760 69.0620 98.1760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9990 142.4100 3.2980 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.0990 142.4100 2.3980 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.3970 142.4100 62.6960 142.7100 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.2980 142.4100 63.5970 142.7100 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3450 0.0000 4.5450 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3450 0.0000 4.5450 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3450 0.0000 4.5450 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3450 0.0000 4.5450 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3450 0.0000 4.5450 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7130 0.0000 5.9130 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7130 0.0000 5.9130 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7130 0.0000 5.9130 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7130 0.0000 5.9130 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7130 0.0000 5.9130 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6090 0.0000 1.8090 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6090 0.0000 1.8090 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6090 0.0000 1.8090 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6090 0.0000 1.8090 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6090 0.0000 1.8090 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9770 0.0000 3.1770 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9770 0.0000 3.1770 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9770 0.0000 3.1770 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9770 0.0000 3.1770 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9770 0.0000 3.1770 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0810 0.0000 7.2810 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0810 0.0000 7.2810 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0810 0.0000 7.2810 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0810 0.0000 7.2810 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0810 0.0000 7.2810 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4490 0.0000 8.6490 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4490 0.0000 8.6490 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4490 0.0000 8.6490 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4490 0.0000 8.6490 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4490 0.0000 8.6490 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8170 0.0000 10.0170 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8170 0.0000 10.0170 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8170 0.0000 10.0170 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8170 0.0000 10.0170 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8170 0.0000 10.0170 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1850 0.0000 11.3850 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1850 0.0000 11.3850 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1850 0.0000 11.3850 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1850 0.0000 11.3850 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1850 0.0000 11.3850 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.9210 0.0000 14.1210 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.9210 0.0000 14.1210 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.9210 0.0000 14.1210 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.9210 0.0000 14.1210 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.9210 0.0000 14.1210 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5530 0.0000 12.7530 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5530 0.0000 12.7530 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5530 0.0000 12.7530 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5530 0.0000 12.7530 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5530 0.0000 12.7530 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.2890 0.0000 15.4890 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.2890 0.0000 15.4890 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.2890 0.0000 15.4890 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.2890 0.0000 15.4890 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.2890 0.0000 15.4890 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.6570 0.0000 16.8570 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.6570 0.0000 16.8570 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.6570 0.0000 16.8570 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.6570 0.0000 16.8570 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.6570 0.0000 16.8570 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.0250 0.0000 18.2250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.0250 0.0000 18.2250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.0250 0.0000 18.2250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.0250 0.0000 18.2250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 19.3930 0.0060 19.5930 0.2060 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.3930 0.0060 19.5930 0.2060 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.3930 0.0060 19.5930 0.2060 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.3930 0.0060 19.5930 0.2060 ;
    END
    PORT
      LAYER M1 ;
        RECT 19.3930 0.0060 19.5930 0.2060 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4970 0.0000 23.6970 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4970 0.0000 23.6970 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4970 0.0000 23.6970 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4970 0.0000 23.6970 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4970 0.0000 23.6970 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0030 0.0000 31.2030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0030 0.0000 31.2030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0030 0.0000 31.2030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0030 0.0000 31.2030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0030 0.0000 31.2030 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442248 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442248 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[6]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.3740 0.0000 32.5740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.3740 0.0000 32.5740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.3760 0.0000 32.5760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.3760 0.0000 32.5760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.3760 0.0000 32.5760 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.354192 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.354192 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[20]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.7420 0.0000 33.9420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.7420 0.0000 33.9420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.7420 0.0000 33.9420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.7420 0.0000 33.9420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.7420 0.0000 33.9420 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[5]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1080 0.0000 35.3080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1080 0.0000 35.3080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1080 0.0000 35.3080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1080 0.0000 35.3080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1080 0.0000 35.3080 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[26]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4750 0.0000 36.6750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4750 0.0000 36.6750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4750 0.0000 36.6750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4750 0.0000 36.6750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4750 0.0000 36.6750 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442248 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442248 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[4]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.8430 0.0000 38.0430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.8430 0.0000 38.0430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.8430 0.0000 38.0430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.8430 0.0000 38.0430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.8430 0.0000 38.0430 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442248 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442248 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[3]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2110 0.0000 39.4110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2110 0.0000 39.4110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2110 0.0000 39.4110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2110 0.0000 39.4110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2110 0.0000 39.4110 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442248 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442248 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[2]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5800 0.0000 40.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5800 0.0000 40.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5800 0.0000 40.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5800 0.0000 40.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5800 0.0000 40.7800 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[1]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.9500 0.0000 42.1500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.9500 0.0000 42.1500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.9510 0.0000 42.1510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.9510 0.0000 42.1510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.9510 0.0000 42.1510 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352457 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352457 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[0]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3160 0.0000 43.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3160 0.0000 43.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3140 0.0000 43.5140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3140 0.0000 43.5140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3140 0.0000 43.5140 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442198 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442198 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[27]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.0480 0.0000 46.2480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.0480 0.0000 46.2480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.0480 0.0000 46.2480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.0480 0.0000 46.2480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.0480 0.0000 46.2480 0.2000 ;
    END
    ANTENNADIFFAREA 18.42974 LAYER M1 ;
    ANTENNADIFFAREA 18.42974 LAYER M2 ;
    ANTENNADIFFAREA 18.42974 LAYER M3 ;
    ANTENNADIFFAREA 18.42974 LAYER M4 ;
    ANTENNADIFFAREA 18.42974 LAYER M5 ;
    ANTENNADIFFAREA 18.42974 LAYER M6 ;
    ANTENNADIFFAREA 18.42974 LAYER M7 ;
    ANTENNADIFFAREA 18.42974 LAYER M8 ;
    ANTENNADIFFAREA 18.42974 LAYER M9 ;
    ANTENNADIFFAREA 18.42974 LAYER MRDL ;
    ANTENNAGATEAREA 2.7159 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 32.76542 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 32.76542 LAYER M1 ;
    ANTENNAGATEAREA 2.7159 LAYER M2 ;
    ANTENNAGATEAREA 2.7159 LAYER M3 ;
    ANTENNAGATEAREA 2.7159 LAYER M4 ;
    ANTENNAGATEAREA 2.7159 LAYER M5 ;
    ANTENNAGATEAREA 2.7159 LAYER M6 ;
    ANTENNAGATEAREA 2.7159 LAYER M7 ;
    ANTENNAGATEAREA 2.7159 LAYER M8 ;
    ANTENNAGATEAREA 2.7159 LAYER M9 ;
    ANTENNAGATEAREA 2.7159 LAYER MRDL ;
  END O[29]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.6880 0.0000 44.8880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.6880 0.0000 44.8880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.6880 0.0000 44.8880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.6880 0.0000 44.8880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.6880 0.0000 44.8880 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352652 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352652 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[28]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4050 0.0000 47.6050 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4050 0.0000 47.6050 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4050 0.0000 47.6050 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4050 0.0000 47.6050 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4050 0.0000 47.6050 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[19]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 9.7900 69.0620 9.9900 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 9.7900 69.0620 9.9900 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 9.7900 69.0620 9.9900 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 9.7900 69.0620 9.9900 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 9.7900 69.0620 9.9900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 87.2230 69.0620 87.4230 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 87.2230 69.0620 87.4230 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 87.2230 69.0620 87.4230 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 87.2230 69.0620 87.4230 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 87.2230 69.0620 87.4230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 90.3480 69.0620 90.5480 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 90.3480 69.0620 90.5480 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 90.3480 69.0620 90.5480 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 90.3480 69.0620 90.5480 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 90.3480 69.0620 90.5480 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 122.8460 69.0620 123.0460 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 122.8460 69.0620 123.0460 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 122.8460 69.0620 123.0460 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 122.8460 69.0620 123.0460 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 122.8460 69.0620 123.0460 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 115.6160 69.0620 115.8160 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 115.6160 69.0620 115.8160 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 115.6160 69.0620 115.8160 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 115.6160 69.0620 115.8160 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 115.6160 69.0620 115.8160 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 114.0260 69.0620 114.2260 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 114.0260 69.0620 114.2260 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 114.0260 69.0620 114.2260 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 114.0260 69.0620 114.2260 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 114.0260 69.0620 114.2260 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.5950 0.0000 14.7950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.5950 0.0000 14.7950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.5950 0.0000 14.7950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.5950 0.0000 14.7950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.5950 0.0000 14.7950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[14]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.0580 0.0000 20.2580 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.0580 0.0000 20.2580 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.0580 0.0000 20.2580 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.0580 0.0000 20.2580 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.0580 0.0000 20.2580 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.443598 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.443598 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[18]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 17.3240 0.0000 17.5240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.3240 0.0000 17.5240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.3240 0.0000 17.5240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 17.3240 0.0000 17.5240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 17.3240 0.0000 17.5240 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[16]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.6920 0.0000 18.8920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.6920 0.0000 18.8920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.6920 0.0000 18.8920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.6920 0.0000 18.8920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.6920 0.0000 18.8920 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[17]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2760 0.0000 2.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2760 0.0000 2.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2760 0.0000 2.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2760 0.0000 2.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2760 0.0000 2.4760 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[30]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.4280 0.0000 21.6280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.4280 0.0000 21.6280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.4280 0.0000 21.6280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.4280 0.0000 21.6280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.4280 0.0000 21.6280 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[21]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.7940 0.0000 22.9940 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.7940 0.0000 22.9940 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.7940 0.0000 22.9940 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.7940 0.0000 22.9940 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.7940 0.0000 22.9940 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442198 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442198 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[7]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.1630 0.0000 24.3630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.1630 0.0000 24.3630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.1630 0.0000 24.3630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.1630 0.0000 24.3630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.1630 0.0000 24.3630 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442248 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442248 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[22]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.5320 0.0000 25.7320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.5320 0.0000 25.7320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.5320 0.0000 25.7320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.5320 0.0000 25.7320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.5320 0.0000 25.7320 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[8]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9000 0.0000 27.1000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9000 0.0000 27.1000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9000 0.0000 27.1000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9000 0.0000 27.1000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9000 0.0000 27.1000 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352312 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352312 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[23]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.2710 0.0000 28.4710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.2710 0.0000 28.4710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.2710 0.0000 28.4710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.2710 0.0000 28.4710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.2710 0.0000 28.4710 0.2000 ;
    END
    ANTENNADIFFAREA 1.582472 LAYER M1 ;
    ANTENNADIFFAREA 1.582472 LAYER M2 ;
    ANTENNADIFFAREA 1.582472 LAYER M3 ;
    ANTENNADIFFAREA 1.582472 LAYER M4 ;
    ANTENNADIFFAREA 1.582472 LAYER M5 ;
    ANTENNADIFFAREA 1.582472 LAYER M6 ;
    ANTENNADIFFAREA 1.582472 LAYER M7 ;
    ANTENNADIFFAREA 1.582472 LAYER M8 ;
    ANTENNADIFFAREA 1.582472 LAYER M9 ;
    ANTENNADIFFAREA 1.582472 LAYER MRDL ;
    ANTENNAGATEAREA 0.2265 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.352457 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.352457 LAYER M1 ;
    ANTENNAGATEAREA 0.2265 LAYER M2 ;
    ANTENNAGATEAREA 0.2265 LAYER M3 ;
    ANTENNAGATEAREA 0.2265 LAYER M4 ;
    ANTENNAGATEAREA 0.2265 LAYER M5 ;
    ANTENNAGATEAREA 0.2265 LAYER M6 ;
    ANTENNAGATEAREA 0.2265 LAYER M7 ;
    ANTENNAGATEAREA 0.2265 LAYER M8 ;
    ANTENNAGATEAREA 0.2265 LAYER M9 ;
    ANTENNAGATEAREA 0.2265 LAYER MRDL ;
  END O[9]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.6350 0.0000 29.8350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.6350 0.0000 29.8350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.6350 0.0000 29.8350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.6350 0.0000 29.8350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.6350 0.0000 29.8350 0.2000 ;
    END
    ANTENNADIFFAREA 1.760972 LAYER M1 ;
    ANTENNADIFFAREA 1.760972 LAYER M2 ;
    ANTENNADIFFAREA 1.760972 LAYER M3 ;
    ANTENNADIFFAREA 1.760972 LAYER M4 ;
    ANTENNADIFFAREA 1.760972 LAYER M5 ;
    ANTENNADIFFAREA 1.760972 LAYER M6 ;
    ANTENNADIFFAREA 1.760972 LAYER M7 ;
    ANTENNADIFFAREA 1.760972 LAYER M8 ;
    ANTENNADIFFAREA 1.760972 LAYER M9 ;
    ANTENNADIFFAREA 1.760972 LAYER MRDL ;
    ANTENNAGATEAREA 0.2445 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 4.442248 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.442248 LAYER M1 ;
    ANTENNAGATEAREA 0.2445 LAYER M2 ;
    ANTENNAGATEAREA 0.2445 LAYER M3 ;
    ANTENNAGATEAREA 0.2445 LAYER M4 ;
    ANTENNAGATEAREA 0.2445 LAYER M5 ;
    ANTENNAGATEAREA 0.2445 LAYER M6 ;
    ANTENNAGATEAREA 0.2445 LAYER M7 ;
    ANTENNAGATEAREA 0.2445 LAYER M8 ;
    ANTENNAGATEAREA 0.2445 LAYER M9 ;
    ANTENNAGATEAREA 0.2445 LAYER MRDL ;
  END O[25]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.9560 0.0000 16.1560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.9560 0.0000 16.1560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.9560 0.0000 16.1560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.9560 0.0000 16.1560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.9560 0.0000 16.1560 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[15]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7480 0.0000 7.9480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7480 0.0000 7.9480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7480 0.0000 7.9480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7480 0.0000 7.9480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7480 0.0000 7.9480 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[10]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.2270 0.0000 13.4270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.2270 0.0000 13.4270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.2270 0.0000 13.4270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.2270 0.0000 13.4270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.2270 0.0000 13.4270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[24]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6440 0.0000 3.8440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6440 0.0000 3.8440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6440 0.0000 3.8440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6440 0.0000 3.8440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6440 0.0000 3.8440 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[31]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.8620 16.4820 69.0620 16.6820 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.8620 16.4820 69.0620 16.6820 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.8620 16.4820 69.0620 16.6820 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.8620 16.4820 69.0620 16.6820 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.8620 16.4820 69.0620 16.6820 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB
  OBS
    LAYER M2 ;
      RECT 0.0000 113.3260 68.1620 116.5160 ;
      RECT 0.0000 107.6960 69.0620 113.3260 ;
      RECT 0.0000 104.5060 68.1620 107.6960 ;
      RECT 0.0000 98.8760 69.0620 104.5060 ;
      RECT 0.0000 97.2760 68.1620 98.8760 ;
      RECT 0.0000 91.2480 69.0620 97.2760 ;
      RECT 0.0000 85.8860 68.1620 91.2480 ;
      RECT 0.0000 17.8940 69.0620 85.8860 ;
      RECT 0.0000 15.7820 68.1620 17.8940 ;
      RECT 0.0000 10.6900 69.0620 15.7820 ;
      RECT 0.0000 9.0900 68.1620 10.6900 ;
      RECT 0.0000 0.9060 69.0620 9.0900 ;
      RECT 0.0000 0.9000 18.6930 0.9060 ;
      RECT 20.2930 0.9000 44.6850 142.7100 ;
      RECT 20.2930 0.9030 69.0620 9.0900 ;
      RECT 20.2930 0.9030 69.0620 0.9060 ;
      RECT 46.2850 0.9000 69.0620 9.0900 ;
      RECT 49.0100 0.0000 69.0620 9.0900 ;
      RECT 0.0000 0.0000 0.9090 0.9000 ;
      RECT 67.5610 88.1230 69.0620 89.6480 ;
      RECT 49.0100 0.0000 69.0620 0.9000 ;
      RECT 20.2930 0.9000 44.6850 0.9030 ;
      RECT 46.2850 0.9000 69.0620 0.9030 ;
      RECT 0.0000 0.9000 18.6930 142.7100 ;
      RECT 0.0000 123.7460 69.0620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 122.1460 68.1620 123.7460 ;
      RECT 0.0000 116.5160 69.0620 122.1460 ;
    LAYER M1 ;
      RECT 68.2620 106.0060 69.0620 106.1960 ;
      RECT 68.2620 114.8260 69.0620 115.0160 ;
      RECT 0.0000 0.0000 1.0090 0.8000 ;
      RECT 67.5610 88.0230 69.0620 89.7480 ;
      RECT 48.9100 0.0000 69.0620 0.8000 ;
      RECT 20.1930 0.8000 44.7850 0.8030 ;
      RECT 46.1850 0.8000 69.0620 0.8030 ;
      RECT 0.0000 0.8000 18.7930 142.7100 ;
      RECT 0.0000 123.6460 69.0620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 0.8060 68.2620 142.7100 ;
      RECT 0.0000 122.2460 68.2620 123.6460 ;
      RECT 0.0000 116.4160 69.0620 122.2460 ;
      RECT 0.0000 113.4260 68.2620 116.4160 ;
      RECT 0.0000 107.5960 69.0620 113.4260 ;
      RECT 0.0000 104.6060 68.2620 107.5960 ;
      RECT 0.0000 98.7760 69.0620 104.6060 ;
      RECT 0.0000 97.3760 68.2620 98.7760 ;
      RECT 0.0000 91.1480 69.0620 97.3760 ;
      RECT 0.0000 85.9860 68.2620 91.1480 ;
      RECT 0.0000 17.7940 69.0620 85.9860 ;
      RECT 0.0000 15.8820 68.2620 17.7940 ;
      RECT 0.0000 10.5900 69.0620 15.8820 ;
      RECT 0.0000 9.1900 68.2620 10.5900 ;
      RECT 0.0000 0.8060 69.0620 9.1900 ;
      RECT 0.0000 0.8000 18.7930 0.8060 ;
      RECT 20.1930 0.8000 44.7850 142.7100 ;
      RECT 20.1930 0.8030 69.0620 9.1900 ;
      RECT 20.1930 0.8030 69.0620 0.8060 ;
      RECT 46.1850 0.8000 69.0620 9.1900 ;
      RECT 48.9100 0.0000 69.0620 9.1900 ;
    LAYER PO ;
      RECT 0.0000 0.0000 69.0620 142.7100 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 69.0620 142.7100 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 69.0620 142.7100 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 69.0620 142.7100 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 69.0620 142.7100 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 69.0620 142.7100 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 0.9090 0.9060 ;
      RECT 0.0000 0.0000 0.9090 0.9000 ;
      RECT 68.3470 141.7100 69.0620 142.7100 ;
      RECT 67.5610 88.1230 69.0620 89.6480 ;
      RECT 49.0100 0.0000 69.0620 0.9000 ;
      RECT 20.2930 0.9000 44.6850 0.9030 ;
      RECT 46.2850 0.9000 69.0620 0.9030 ;
      RECT 0.0000 0.9000 18.6930 141.7100 ;
      RECT 0.0000 123.7460 69.0620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 0.9060 68.1620 141.7100 ;
      RECT 0.0000 122.1460 68.1620 123.7460 ;
      RECT 0.0000 116.5160 69.0620 122.1460 ;
      RECT 0.0000 113.3260 68.1620 116.5160 ;
      RECT 0.0000 107.6960 69.0620 113.3260 ;
      RECT 0.0000 104.5060 68.1620 107.6960 ;
      RECT 0.0000 98.8760 69.0620 104.5060 ;
      RECT 0.0000 97.2760 68.1620 98.8760 ;
      RECT 0.0000 91.2480 69.0620 97.2760 ;
      RECT 0.0000 85.8860 68.1620 91.2480 ;
      RECT 0.0000 17.8940 69.0620 85.8860 ;
      RECT 0.0000 15.7820 68.1620 17.8940 ;
      RECT 0.0000 10.6900 69.0620 15.7820 ;
      RECT 0.0000 9.0900 68.1620 10.6900 ;
      RECT 0.0000 0.9060 69.0620 9.0900 ;
      RECT 0.0000 0.9000 18.6930 0.9060 ;
      RECT 20.2930 0.9000 44.6850 141.7100 ;
      RECT 20.2930 0.9030 69.0620 9.0900 ;
      RECT 20.2930 0.9030 69.0620 0.9060 ;
      RECT 46.2850 0.9000 69.0620 9.0900 ;
      RECT 49.0100 0.0000 69.0620 9.0900 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9090 0.9060 ;
      RECT 0.0000 0.0000 0.9090 0.9000 ;
      RECT 67.5610 88.1230 69.0620 89.6480 ;
      RECT 49.0100 0.0000 69.0620 0.9000 ;
      RECT 20.2930 0.9000 44.6850 0.9030 ;
      RECT 46.2850 0.9000 69.0620 0.9030 ;
      RECT 0.0000 0.9000 18.6930 142.7100 ;
      RECT 0.0000 123.7460 69.0620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 122.1460 68.1620 123.7460 ;
      RECT 0.0000 116.5160 69.0620 122.1460 ;
      RECT 0.0000 113.3260 68.1620 116.5160 ;
      RECT 0.0000 107.6960 69.0620 113.3260 ;
      RECT 0.0000 104.5060 68.1620 107.6960 ;
      RECT 0.0000 98.8760 69.0620 104.5060 ;
      RECT 0.0000 97.2760 68.1620 98.8760 ;
      RECT 0.0000 91.2480 69.0620 97.2760 ;
      RECT 0.0000 85.8860 68.1620 91.2480 ;
      RECT 0.0000 17.8940 69.0620 85.8860 ;
      RECT 0.0000 15.7820 68.1620 17.8940 ;
      RECT 0.0000 10.6900 69.0620 15.7820 ;
      RECT 0.0000 9.0900 68.1620 10.6900 ;
      RECT 0.0000 0.9060 69.0620 9.0900 ;
      RECT 0.0000 0.9000 18.6930 0.9060 ;
      RECT 20.2930 0.9000 44.6850 142.7100 ;
      RECT 20.2930 0.9030 69.0620 9.0900 ;
      RECT 20.2930 0.9030 69.0620 0.9060 ;
      RECT 46.2850 0.9000 69.0620 9.0900 ;
      RECT 49.0100 0.0000 69.0620 9.0900 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9090 0.9060 ;
      RECT 0.0000 0.0000 0.9090 0.9000 ;
      RECT 67.5610 88.1230 69.0620 89.6480 ;
      RECT 49.0100 0.0000 69.0620 0.9000 ;
      RECT 20.2930 0.9000 44.6850 0.9030 ;
      RECT 46.2850 0.9000 69.0620 0.9030 ;
      RECT 0.0000 0.9000 18.6930 142.7100 ;
      RECT 0.0000 123.7460 69.0620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 0.9060 68.1620 142.7100 ;
      RECT 0.0000 122.1460 68.1620 123.7460 ;
      RECT 0.0000 116.5160 69.0620 122.1460 ;
      RECT 0.0000 113.3260 68.1620 116.5160 ;
      RECT 0.0000 107.6960 69.0620 113.3260 ;
      RECT 0.0000 104.5060 68.1620 107.6960 ;
      RECT 0.0000 98.8760 69.0620 104.5060 ;
      RECT 0.0000 97.2760 68.1620 98.8760 ;
      RECT 0.0000 91.2480 69.0620 97.2760 ;
      RECT 0.0000 85.8860 68.1620 91.2480 ;
      RECT 0.0000 17.8940 69.0620 85.8860 ;
      RECT 0.0000 15.7820 68.1620 17.8940 ;
      RECT 0.0000 10.6900 69.0620 15.7820 ;
      RECT 0.0000 9.0900 68.1620 10.6900 ;
      RECT 0.0000 0.9060 69.0620 9.0900 ;
      RECT 0.0000 0.9000 18.6930 0.9060 ;
      RECT 20.2930 0.9000 44.6850 142.7100 ;
      RECT 20.2930 0.9030 69.0620 9.0900 ;
      RECT 20.2930 0.9030 69.0620 0.9060 ;
      RECT 46.2850 0.9000 69.0620 9.0900 ;
      RECT 49.0100 0.0000 69.0620 9.0900 ;
  END
END SRAMLP1RW64x34

MACRO SRAMLP1RW64x128
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 197.522 BY 140.744 ;
  SYMMETRY X Y R90 ;

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[29]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[26]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[25]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[26]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[27]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[27]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[43]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[42]

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[44]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[41]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[41]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[40]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[40]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[42]

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[38]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[39]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[37]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[39]

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[38]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[37]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[36]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[35]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[36]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[34]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 98.7070 197.5220 98.9070 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 98.7070 197.5220 98.9070 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 98.7070 197.5220 98.9070 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 98.7070 197.5220 98.9070 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 98.7070 197.5220 98.9070 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[5]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 176.7010 0.0000 176.9010 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.7010 0.0000 176.9010 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.7010 0.0000 176.9010 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 176.7010 0.0000 176.9010 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 176.7010 0.0000 176.9010 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END OEB

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 17.2900 197.5220 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 17.2900 197.5220 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 17.2900 197.5220 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 17.2900 197.5220 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 17.2900 197.5220 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CE

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[45]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[43]

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 107.6230 197.5220 107.8230 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 107.6230 197.5220 107.8230 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 107.6230 197.5220 107.8230 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 107.6230 197.5220 107.8230 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 107.6230 197.5220 107.8230 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[3]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 116.4550 197.5220 116.6550 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 116.4550 197.5220 116.6550 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 116.4550 197.5220 116.6550 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 116.4550 197.5220 116.6550 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 116.4550 197.5220 116.6550 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[1]

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 123.6850 197.5220 123.8850 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 123.6850 197.5220 123.8850 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 123.6850 197.5220 123.8850 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 123.6850 197.5220 123.8850 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 123.6850 197.5220 123.8850 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[0]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 106.0450 197.5220 106.2450 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 106.0450 197.5220 106.2450 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 106.0450 197.5220 106.2450 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 106.0450 197.5220 106.2450 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 106.0450 197.5220 106.2450 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[4]

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 114.8650 197.5220 115.0650 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 114.8650 197.5220 115.0650 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 114.8650 197.5220 115.0650 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 114.8650 197.5220 115.0650 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 114.8650 197.5220 115.0650 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END A[2]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 3.1610 140.4440 3.4620 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.2620 140.4440 2.5610 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.9610 140.4440 194.2600 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.8610 140.4440 195.1610 140.7440 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 1.8110 140.4440 2.1110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.7130 140.4440 3.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.6130 140.4440 3.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.9120 140.4440 1.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.1120 140.4440 8.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.2120 140.4440 7.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.4120 140.4440 5.7130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.3120 140.4440 6.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.5130 140.4440 4.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.6120 140.4440 12.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.0130 140.4440 9.3130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.8130 140.4440 11.1140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.7120 140.4440 12.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.9120 140.4440 10.2110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.1120 140.4440 17.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.5130 140.4440 13.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.4120 140.4440 14.7110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.2120 140.4440 16.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.0130 140.4440 18.3130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.3130 140.4440 15.6140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.6120 140.4440 21.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.9120 140.4440 19.2110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.8130 140.4440 20.1140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.5130 140.4440 22.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.7120 140.4440 21.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.9120 140.4440 28.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.0120 140.4440 27.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.2120 140.4440 25.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.3120 140.4440 24.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.4120 140.4440 23.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.1130 140.4440 26.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.4110 140.4440 32.7110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.5120 140.4440 31.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.6120 140.4440 30.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.8120 140.4440 29.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.7130 140.4440 30.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.2110 140.4440 34.5110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.1130 140.4440 35.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.0130 140.4440 36.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.9130 140.4440 37.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.3120 140.4440 33.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.5120 140.4440 40.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.6120 140.4440 39.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.4130 140.4440 41.7130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.8120 140.4440 38.1130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.3120 140.4440 42.6110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.7120 140.4440 39.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.0120 140.4440 45.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.9130 140.4440 46.2130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.8120 140.4440 47.1110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.2130 140.4440 43.5140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.1120 140.4440 44.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.5120 140.4440 49.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.6120 140.4440 48.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.3120 140.4440 51.6110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.4130 140.4440 50.7130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.7130 140.4440 48.0140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.7120 140.4440 57.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.8120 140.4440 56.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.0120 140.4440 54.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.2130 140.4440 52.5140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.9130 140.4440 55.2130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.1120 140.4440 53.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.2120 140.4440 61.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.3120 140.4440 60.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.4120 140.4440 59.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.6120 140.4440 57.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.5130 140.4440 58.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.8110 140.4440 65.1110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.9120 140.4440 64.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.0120 140.4440 63.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.7120 140.4440 66.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.1130 140.4440 62.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.2120 140.4440 70.5130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.6110 140.4440 66.9110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.5130 140.4440 67.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.1120 140.4440 71.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.4130 140.4440 68.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.3130 140.4440 69.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.9120 140.4440 73.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.0120 140.4440 72.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.8130 140.4440 74.1130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.6130 140.4440 75.9140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.7120 140.4440 75.0110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.4120 140.4440 77.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.3130 140.4440 78.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.2120 140.4440 79.5110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.5120 140.4440 76.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.1130 140.4440 80.4140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.9120 140.4440 82.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.0120 140.4440 81.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.7120 140.4440 84.0110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.8130 140.4440 83.1130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.6130 140.4440 84.9140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.5120 140.4440 85.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.0120 140.4440 90.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.1120 140.4440 89.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.2120 140.4440 88.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.4120 140.4440 86.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.3130 140.4440 87.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.6120 140.4440 93.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.7120 140.4440 93.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.8120 140.4440 92.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.5130 140.4440 94.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.9130 140.4440 91.2130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.0110 140.4440 99.3110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.2110 140.4440 97.5110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.3120 140.4440 96.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.4120 140.4440 95.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.9130 140.4440 100.2130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.1120 140.4440 98.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.4120 140.4440 104.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.6120 140.4440 102.9130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.5120 140.4440 103.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.8130 140.4440 101.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.7130 140.4440 102.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.3120 140.4440 105.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.8120 140.4440 110.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.2130 140.4440 106.5130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.0130 140.4440 108.3140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.9120 140.4440 109.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.1120 140.4440 107.4110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.3120 140.4440 114.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.7130 140.4440 111.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.6120 140.4440 111.9110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.4120 140.4440 113.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.5130 140.4440 112.8140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.8120 140.4440 119.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.1120 140.4440 116.4110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.2130 140.4440 115.5130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.0130 140.4440 117.3140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.9120 140.4440 118.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.2120 140.4440 124.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.4120 140.4440 122.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.5120 140.4440 121.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.6120 140.4440 120.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.3130 140.4440 123.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.7130 140.4440 120.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.7120 140.4440 129.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.8120 140.4440 128.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.0120 140.4440 126.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.1120 140.4440 125.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.9130 140.4440 127.2130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.3130 140.4440 132.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.2130 140.4440 133.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.5120 140.4440 130.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.4110 140.4440 131.7110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.6110 140.4440 129.9110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.7120 140.4440 138.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.8120 140.4440 137.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.6130 140.4440 138.9130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.0120 140.4440 135.3130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.9120 140.4440 136.2130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.1130 140.4440 134.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.2120 140.4440 142.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.1130 140.4440 143.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.4130 140.4440 140.7140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.3120 140.4440 141.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.5120 140.4440 139.8110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.0120 140.4440 144.3110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.8120 140.4440 146.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.6130 140.4440 147.9130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.7120 140.4440 147.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.9130 140.4440 145.2140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.5120 140.4440 148.8110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.4130 140.4440 149.7140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.1130 140.4440 152.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.3120 140.4440 150.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.0120 140.4440 153.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.2120 140.4440 151.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.7130 140.4440 156.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.5120 140.4440 157.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.6120 140.4440 156.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.8120 140.4440 155.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.9120 140.4440 154.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.3130 140.4440 159.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.0110 140.4440 162.3110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.1120 140.4440 161.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.2120 140.4440 160.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.4120 140.4440 158.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.4120 140.4440 167.7130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.7130 140.4440 165.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.6130 140.4440 165.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.5130 140.4440 166.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.9120 140.4440 163.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 163.8110 140.4440 164.1110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.1120 140.4440 170.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.2120 140.4440 169.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.0130 140.4440 171.3130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.9120 140.4440 172.2110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.3120 140.4440 168.6130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 174.6120 140.4440 174.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.5130 140.4440 175.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.4120 140.4440 176.7110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.8130 140.4440 173.1140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.7120 140.4440 174.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.2120 140.4440 178.5120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.9120 140.4440 181.2110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.0130 140.4440 180.3130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.8130 140.4440 182.1140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.1120 140.4440 179.4120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.3130 140.4440 177.6140 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.5130 140.4440 184.8130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.7120 140.4440 183.0120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.3120 140.4440 186.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 185.4120 140.4440 185.7120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.6120 140.4440 183.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.1130 140.4440 188.4130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.8120 140.4440 191.1120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.9120 140.4440 190.2120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.0120 140.4440 189.3120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.6120 140.4440 192.9120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.5120 140.4440 193.8120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.4110 140.4440 194.7110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.2110 140.4440 196.5110 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 191.7130 140.4440 192.0130 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 195.3120 140.4440 195.6120 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 187.2120 140.4440 187.5120 140.7440 ;
    END
  END VSS

  PIN I[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.1110 0.0000 74.3110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.1110 0.0000 74.3110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.1110 0.0000 74.3110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.1110 0.0000 74.3110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.1110 0.0000 74.3110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[53]

  PIN O[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 74.7960 0.0000 74.9960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.7960 0.0000 74.9960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.7960 0.0000 74.9960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 74.7960 0.0000 74.9960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 74.7960 0.0000 74.9960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[53]

  PIN I[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 75.4790 0.0000 75.6790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.4790 0.0000 75.6790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.4790 0.0000 75.6790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 75.4790 0.0000 75.6790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 75.4790 0.0000 75.6790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[54]

  PIN O[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.1640 0.0000 76.3640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.1640 0.0000 76.3640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.1640 0.0000 76.3640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.1640 0.0000 76.3640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.1640 0.0000 76.3640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[54]

  PIN I[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 76.8470 0.0000 77.0470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.8470 0.0000 77.0470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.8470 0.0000 77.0470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 76.8470 0.0000 77.0470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 76.8470 0.0000 77.0470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[55]

  PIN O[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 77.5320 0.0000 77.7320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.5320 0.0000 77.7320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.5320 0.0000 77.7320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 77.5320 0.0000 77.7320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 77.5320 0.0000 77.7320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[55]

  PIN I[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.2150 0.0000 78.4150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.2150 0.0000 78.4150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.2150 0.0000 78.4150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.2150 0.0000 78.4150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.2150 0.0000 78.4150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[56]

  PIN O[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 78.9000 0.0000 79.1000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.9000 0.0000 79.1000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.9000 0.0000 79.1000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 78.9000 0.0000 79.1000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 78.9000 0.0000 79.1000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[56]

  PIN I[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 79.5830 0.0000 79.7830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.5830 0.0000 79.7830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.5830 0.0000 79.7830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 79.5830 0.0000 79.7830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 79.5830 0.0000 79.7830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[57]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[7]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[2]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[4]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[4]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[3]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[5]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN I[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.2710 0.0000 67.4710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[48]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[0]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9750 0.0010 3.1750 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9750 0.0010 3.1750 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[1]

  PIN I[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5350 0.0000 64.7350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[46]

  PIN O[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.2200 0.0000 65.4200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[46]

  PIN I[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 65.9030 0.0010 66.1030 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.9030 0.0010 66.1030 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 65.9030 0.0000 66.1030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[47]

  PIN O[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 66.5880 0.0000 66.7880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[47]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3280 133.6430 197.5220 133.8430 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3280 133.6430 197.5220 133.8430 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3280 133.6430 197.5220 133.8430 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3280 133.6430 197.5220 133.8430 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3280 133.6430 197.5220 133.8430 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END LS

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[14]

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[12]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[13]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[11]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[10]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[9]

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[8]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[6]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[24]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[22]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[23]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[18]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[19]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[21]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[20]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[17]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[16]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[15]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[33]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[32]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[31]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[30]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[29]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[28]

  PIN O[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 122.6760 0.0000 122.8760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.6760 0.0000 122.8760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.6760 0.0000 122.8760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 122.6760 0.0000 122.8760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 122.6760 0.0000 122.8760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[88]

  PIN I[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 123.3590 0.0000 123.5590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.3590 0.0000 123.5590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.3590 0.0000 123.5590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 123.3590 0.0000 123.5590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 123.3590 0.0000 123.5590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[89]

  PIN O[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 124.0440 0.0000 124.2440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.0440 0.0000 124.2440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.0440 0.0000 124.2440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 124.0440 0.0000 124.2440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.0440 0.0000 124.2440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[89]

  PIN I[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 124.7270 0.0000 124.9270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.7270 0.0000 124.9270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.7270 0.0000 124.9270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 124.7270 0.0000 124.9270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 124.7270 0.0000 124.9270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[90]

  PIN O[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 125.4120 0.0000 125.6120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.4120 0.0000 125.6120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.4120 0.0000 125.6120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 125.4120 0.0000 125.6120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 125.4120 0.0000 125.6120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[90]

  PIN I[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 126.0950 0.0000 126.2950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.0950 0.0000 126.2950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.0950 0.0000 126.2950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 126.0950 0.0000 126.2950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 126.0950 0.0000 126.2950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[91]

  PIN O[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 126.7800 0.0000 126.9800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.7800 0.0000 126.9800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.7800 0.0000 126.9800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 126.7800 0.0000 126.9800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 126.7800 0.0000 126.9800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[91]

  PIN I[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 127.4630 0.0000 127.6630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.4630 0.0000 127.6630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.4630 0.0000 127.6630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 127.4630 0.0000 127.6630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 127.4630 0.0000 127.6630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[92]

  PIN O[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 128.1480 0.0000 128.3480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.1480 0.0000 128.3480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.1480 0.0000 128.3480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 128.1480 0.0000 128.3480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 128.1480 0.0000 128.3480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[92]

  PIN I[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 128.8310 0.0010 129.0310 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.8310 0.0010 129.0310 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.8310 0.0000 129.0310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 128.8310 0.0000 129.0310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 128.8310 0.0000 129.0310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[93]

  PIN O[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 129.5160 0.0000 129.7160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.5160 0.0000 129.7160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.5160 0.0000 129.7160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 129.5160 0.0000 129.7160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 129.5160 0.0000 129.7160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[93]

  PIN O[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 136.3560 0.0000 136.5560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.3560 0.0000 136.5560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.3560 0.0000 136.5560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 136.3560 0.0000 136.5560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 136.3560 0.0000 136.5560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[98]

  PIN O[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 130.8840 0.0000 131.0840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.8840 0.0000 131.0840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.8840 0.0000 131.0840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 130.8840 0.0000 131.0840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 130.8840 0.0000 131.0840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[94]

  PIN O[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.2600 0.0000 106.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.2600 0.0000 106.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.2600 0.0000 106.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.2600 0.0000 106.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.2600 0.0000 106.4600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[76]

  PIN I[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 106.9430 0.0000 107.1430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.9430 0.0000 107.1430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.9430 0.0000 107.1430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 106.9430 0.0000 107.1430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 106.9430 0.0000 107.1430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[77]

  PIN O[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 107.6280 0.0000 107.8280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.6280 0.0000 107.8280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.6280 0.0000 107.8280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 107.6280 0.0000 107.8280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 107.6280 0.0000 107.8280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[77]

  PIN I[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.3110 0.0000 108.5110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.3110 0.0000 108.5110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.3110 0.0000 108.5110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.3110 0.0000 108.5110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.3110 0.0000 108.5110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[78]

  PIN O[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 108.9960 0.0000 109.1960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.9960 0.0000 109.1960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.9960 0.0000 109.1960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 108.9960 0.0000 109.1960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 108.9960 0.0000 109.1960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[78]

  PIN I[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 109.6790 0.0000 109.8790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.6790 0.0000 109.8790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.6790 0.0000 109.8790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 109.6790 0.0000 109.8790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 109.6790 0.0000 109.8790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[79]

  PIN O[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 110.3640 0.0000 110.5640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.3640 0.0000 110.5640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.3640 0.0000 110.5640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 110.3640 0.0000 110.5640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 110.3640 0.0000 110.5640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[79]

  PIN I[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.0470 0.0000 111.2470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.0470 0.0000 111.2470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.0470 0.0000 111.2470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.0470 0.0000 111.2470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.0470 0.0000 111.2470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[80]

  PIN O[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 111.7320 0.0000 111.9320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.7320 0.0000 111.9320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.7320 0.0000 111.9320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 111.7320 0.0000 111.9320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 111.7320 0.0000 111.9320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[80]

  PIN I[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 112.4150 0.0000 112.6150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.4150 0.0000 112.6150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.4150 0.0000 112.6150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 112.4150 0.0000 112.6150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 112.4150 0.0000 112.6150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[81]

  PIN O[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 113.1000 0.0000 113.3000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.1000 0.0000 113.3000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.1000 0.0000 113.3000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 113.1000 0.0000 113.3000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.1000 0.0000 113.3000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[81]

  PIN I[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 113.7830 0.0000 113.9830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.7830 0.0000 113.9830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.7830 0.0000 113.9830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 113.7830 0.0000 113.9830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 113.7830 0.0000 113.9830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[82]

  PIN O[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 114.4680 0.0000 114.6680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.4680 0.0000 114.6680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.4680 0.0000 114.6680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 114.4680 0.0000 114.6680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 114.4680 0.0000 114.6680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[82]

  PIN I[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 115.1510 0.0000 115.3510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.1510 0.0000 115.3510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.1510 0.0000 115.3510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.1510 0.0000 115.3510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.1510 0.0000 115.3510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[83]

  PIN O[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 115.8360 0.0000 116.0360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.8360 0.0000 116.0360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.8360 0.0000 116.0360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 115.8360 0.0000 116.0360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 115.8360 0.0000 116.0360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[83]

  PIN I[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 116.5190 0.0000 116.7190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.5190 0.0000 116.7190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.5190 0.0000 116.7190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 116.5190 0.0000 116.7190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 116.5190 0.0000 116.7190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[84]

  PIN O[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 117.2040 0.0000 117.4040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.2040 0.0000 117.4040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.2040 0.0000 117.4040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 117.2040 0.0000 117.4040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.2040 0.0000 117.4040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[84]

  PIN I[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 117.8870 0.0000 118.0870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.8870 0.0000 118.0870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.8870 0.0000 118.0870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 117.8870 0.0000 118.0870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 117.8870 0.0000 118.0870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[85]

  PIN I[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.2630 0.0000 93.4630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.2630 0.0000 93.4630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.2630 0.0000 93.4630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.2630 0.0000 93.4630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.2630 0.0000 93.4630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[67]

  PIN O[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.9480 0.0000 94.1480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.9480 0.0000 94.1480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.9480 0.0000 94.1480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.9480 0.0000 94.1480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.9480 0.0000 94.1480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[67]

  PIN I[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 94.6310 0.0000 94.8310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.6310 0.0000 94.8310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.6310 0.0000 94.8310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 94.6310 0.0000 94.8310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 94.6310 0.0000 94.8310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[68]

  PIN O[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.3160 0.0000 95.5160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.3160 0.0000 95.5160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.3160 0.0000 95.5160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.3160 0.0000 95.5160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.3160 0.0000 95.5160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[68]

  PIN I[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 95.9990 0.0000 96.1990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.9990 0.0000 96.1990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.9990 0.0000 96.1990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 95.9990 0.0000 96.1990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 95.9990 0.0000 96.1990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[69]

  PIN O[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 96.6840 0.0000 96.8840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.6840 0.0000 96.8840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.6840 0.0000 96.8840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 96.6840 0.0000 96.8840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 96.6840 0.0000 96.8840 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[69]

  PIN I[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 97.3670 0.0000 97.5670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.3670 0.0000 97.5670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.3670 0.0000 97.5670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 97.3670 0.0000 97.5670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 97.3670 0.0000 97.5670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[70]

  PIN O[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.0520 0.0000 98.2520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.0520 0.0000 98.2520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.0520 0.0000 98.2520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.0520 0.0000 98.2520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.0520 0.0000 98.2520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[70]

  PIN I[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 98.7350 0.0000 98.9350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.7350 0.0000 98.9350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.7350 0.0000 98.9350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 98.7350 0.0000 98.9350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 98.7350 0.0000 98.9350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[71]

  PIN O[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 99.4200 0.0000 99.6200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.4200 0.0000 99.6200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.4200 0.0000 99.6200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 99.4200 0.0000 99.6200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 99.4200 0.0000 99.6200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[71]

  PIN I[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.1030 0.0000 100.3030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.1030 0.0000 100.3030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.1030 0.0000 100.3030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.1030 0.0000 100.3030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.1030 0.0000 100.3030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[72]

  PIN O[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 100.7880 0.0000 100.9880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.7880 0.0000 100.9880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.7880 0.0000 100.9880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 100.7880 0.0000 100.9880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 100.7880 0.0000 100.9880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[72]

  PIN I[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 101.4710 0.0000 101.6710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.4710 0.0000 101.6710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.4710 0.0000 101.6710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 101.4710 0.0000 101.6710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 101.4710 0.0000 101.6710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[73]

  PIN O[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.1560 0.0000 102.3560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.1560 0.0000 102.3560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.1560 0.0000 102.3560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.1560 0.0000 102.3560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.1560 0.0000 102.3560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[73]

  PIN I[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 102.8390 0.0000 103.0390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.8390 0.0000 103.0390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.8390 0.0000 103.0390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 102.8390 0.0000 103.0390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 102.8390 0.0000 103.0390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[74]

  PIN O[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 103.5240 0.0000 103.7240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.5240 0.0000 103.7240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.5240 0.0000 103.7240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 103.5240 0.0000 103.7240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 103.5240 0.0000 103.7240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[74]

  PIN I[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.2070 0.0000 104.4070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.2070 0.0000 104.4070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.2070 0.0000 104.4070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.2070 0.0000 104.4070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.2070 0.0000 104.4070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[75]

  PIN O[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 104.8920 0.0000 105.0920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.8920 0.0000 105.0920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.8920 0.0000 105.0920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 104.8920 0.0000 105.0920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 104.8920 0.0000 105.0920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[75]

  PIN I[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 105.5750 0.0000 105.7750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.5750 0.0000 105.7750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.5750 0.0000 105.7750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 105.5750 0.0000 105.7750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 105.5750 0.0000 105.7750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[76]

  PIN O[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.2680 0.0000 80.4680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.2680 0.0000 80.4680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.2680 0.0000 80.4680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.2680 0.0000 80.4680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.2680 0.0000 80.4680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[57]

  PIN I[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 80.9510 0.0000 81.1510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.9510 0.0000 81.1510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.9510 0.0000 81.1510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 80.9510 0.0000 81.1510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 80.9510 0.0000 81.1510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[58]

  PIN O[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 81.6360 0.0000 81.8360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.6360 0.0000 81.8360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.6360 0.0000 81.8360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 81.6360 0.0000 81.8360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 81.6360 0.0000 81.8360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[58]

  PIN I[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.6870 0.0000 83.8870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.6870 0.0000 83.8870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.6870 0.0000 83.8870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.6870 0.0000 83.8870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.6870 0.0000 83.8870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[60]

  PIN O[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 84.3720 0.0000 84.5720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.3720 0.0000 84.5720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.3720 0.0000 84.5720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 84.3720 0.0000 84.5720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 84.3720 0.0000 84.5720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[60]

  PIN I[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 82.3190 0.0000 82.5190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.3190 0.0000 82.5190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.3190 0.0000 82.5190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 82.3190 0.0000 82.5190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 82.3190 0.0000 82.5190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[59]

  PIN O[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 83.0040 0.0000 83.2040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.0040 0.0000 83.2040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.0040 0.0000 83.2040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 83.0040 0.0000 83.2040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 83.0040 0.0000 83.2040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[59]

  PIN I[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.0550 0.0000 85.2550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.0550 0.0000 85.2550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.0550 0.0000 85.2550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.0550 0.0000 85.2550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.0550 0.0000 85.2550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[61]

  PIN O[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 85.7400 0.0000 85.9400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.7400 0.0000 85.9400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.7400 0.0000 85.9400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 85.7400 0.0000 85.9400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 85.7400 0.0000 85.9400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[61]

  PIN I[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 86.4230 0.0000 86.6230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.4230 0.0000 86.6230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.4230 0.0000 86.6230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 86.4230 0.0000 86.6230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 86.4230 0.0000 86.6230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[62]

  PIN O[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.1080 0.0000 87.3080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.1080 0.0000 87.3080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.1080 0.0000 87.3080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.1080 0.0000 87.3080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.1080 0.0000 87.3080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[62]

  PIN I[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 87.7910 0.0000 87.9910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.7910 0.0000 87.9910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.7910 0.0000 87.9910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 87.7910 0.0000 87.9910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 87.7910 0.0000 87.9910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[63]

  PIN O[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 88.4760 0.0000 88.6760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.4760 0.0000 88.6760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.4760 0.0000 88.6760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 88.4760 0.0000 88.6760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 88.4760 0.0000 88.6760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[63]

  PIN I[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.1590 0.0000 89.3590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.1590 0.0000 89.3590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.1590 0.0000 89.3590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.1590 0.0000 89.3590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.1590 0.0000 89.3590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[64]

  PIN O[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 89.8440 0.0000 90.0440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.8440 0.0000 90.0440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.8440 0.0000 90.0440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 89.8440 0.0000 90.0440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 89.8440 0.0000 90.0440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[64]

  PIN I[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 90.5270 0.0000 90.7270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.5270 0.0000 90.7270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.5270 0.0000 90.7270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 90.5270 0.0000 90.7270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 90.5270 0.0000 90.7270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[65]

  PIN O[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.2120 0.0000 91.4120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.2120 0.0000 91.4120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.2120 0.0000 91.4120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.2120 0.0000 91.4120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.2120 0.0000 91.4120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[65]

  PIN I[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 91.8950 0.0000 92.0950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.8950 0.0000 92.0950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.8950 0.0000 92.0950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 91.8950 0.0000 92.0950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 91.8950 0.0000 92.0950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[66]

  PIN O[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 92.5800 0.0000 92.7800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.5800 0.0000 92.7800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.5800 0.0000 92.7800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 92.5800 0.0000 92.7800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 92.5800 0.0000 92.7800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[66]

  PIN O[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 67.9560 0.0000 68.1560 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[48]

  PIN I[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 68.6390 0.0000 68.8390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[49]

  PIN O[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 69.3240 0.0000 69.5240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[49]

  PIN I[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.0070 0.0000 70.2070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.0070 0.0000 70.2070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.0070 0.0000 70.2070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.0070 0.0000 70.2070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.0070 0.0000 70.2070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[50]

  PIN O[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 70.6920 0.0000 70.8920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.6920 0.0000 70.8920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.6920 0.0000 70.8920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 70.6920 0.0000 70.8920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 70.6920 0.0000 70.8920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[50]

  PIN I[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 71.3750 0.0000 71.5750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.3750 0.0000 71.5750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.3750 0.0000 71.5750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 71.3750 0.0000 71.5750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 71.3750 0.0000 71.5750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[51]

  PIN O[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.0600 0.0000 72.2600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.0600 0.0000 72.2600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.0600 0.0000 72.2600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.0600 0.0000 72.2600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.0600 0.0000 72.2600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[51]

  PIN I[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 72.7430 0.0000 72.9430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.7430 0.0000 72.9430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.7430 0.0000 72.9430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 72.7430 0.0000 72.9430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 72.7430 0.0000 72.9430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[52]

  PIN O[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 73.4280 0.0000 73.6280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.4280 0.0000 73.6280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.4280 0.0000 73.6280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 73.4280 0.0000 73.6280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 73.4280 0.0000 73.6280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[52]

  PIN I[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 169.8710 0.0000 170.0710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.8710 0.0000 170.0710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.8710 0.0000 170.0710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 169.8710 0.0000 170.0710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 169.8710 0.0000 170.0710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[123]

  PIN O[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 170.5560 0.0000 170.7560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 170.5560 0.0000 170.7560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 170.5560 0.0000 170.7560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 170.5560 0.0000 170.7560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 170.5560 0.0000 170.7560 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[123]

  PIN I[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 171.2390 0.0000 171.4390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.2390 0.0000 171.4390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.2390 0.0000 171.4390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 171.2390 0.0000 171.4390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 171.2390 0.0000 171.4390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[124]

  PIN O[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 171.9240 0.0000 172.1240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.9240 0.0000 172.1240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.9240 0.0000 172.1240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 171.9240 0.0000 172.1240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 171.9240 0.0000 172.1240 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[124]

  PIN I[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 172.6070 0.0000 172.8070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 172.6070 0.0000 172.8070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 172.6070 0.0000 172.8070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 172.6070 0.0000 172.8070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 172.6070 0.0000 172.8070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[125]

  PIN O[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 173.2920 0.0000 173.4920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.2920 0.0000 173.4920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.2920 0.0000 173.4920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 173.2920 0.0000 173.4920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 173.2920 0.0000 173.4920 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[125]

  PIN I[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 173.9750 0.0000 174.1750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.9750 0.0000 174.1750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.9750 0.0000 174.1750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 173.9750 0.0000 174.1750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 173.9750 0.0000 174.1750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[126]

  PIN O[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 174.6600 0.0000 174.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 174.6600 0.0000 174.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 174.6600 0.0000 174.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 174.6600 0.0000 174.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 174.6600 0.0000 174.8600 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[126]

  PIN I[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 175.3430 0.0000 175.5430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.3430 0.0000 175.5430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.3430 0.0000 175.5430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 175.3430 0.0000 175.5430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 175.3430 0.0000 175.5430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[127]

  PIN O[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 176.0280 0.0000 176.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.0280 0.0000 176.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.0280 0.0000 176.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 176.0280 0.0000 176.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 176.0280 0.0000 176.2280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[127]

  PIN VDDL
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.0610 140.4440 4.3620 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.9620 140.4440 5.2620 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.1610 140.4440 192.4600 140.7440 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.0610 140.4440 193.3600 140.7440 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END VDDL

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3280 130.3910 197.5220 130.5910 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3280 130.3910 197.5220 130.5910 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3280 130.3910 197.5220 130.5910 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3280 130.3910 197.5220 130.5910 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3280 130.3910 197.5220 130.5910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END DS

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3280 130.0480 197.5220 130.2480 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3280 130.0480 197.5220 130.2480 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3280 130.0480 197.5220 130.2480 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3280 130.0480 197.5220 130.2480 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3280 130.0480 197.5220 130.2480 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END SD

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3210 9.8200 197.5210 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3210 9.8200 197.5210 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3210 9.8200 197.5210 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3210 9.8200 197.5210 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3210 9.8200 197.5210 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END WEB

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 197.3220 16.8280 197.5220 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.3220 16.8280 197.5220 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.3220 16.8280 197.5220 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 197.3220 16.8280 197.5220 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 197.3220 16.8280 197.5220 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END CSB

  PIN O[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 156.8760 0.0000 157.0760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.8760 0.0000 157.0760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.8760 0.0000 157.0760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 156.8760 0.0000 157.0760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 156.8760 0.0000 157.0760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[113]

  PIN I[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 157.5590 0.0000 157.7590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 157.5590 0.0000 157.7590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 157.5590 0.0000 157.7590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 157.5590 0.0000 157.7590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 157.5590 0.0000 157.7590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[114]

  PIN O[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.2440 0.0000 158.4440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.2440 0.0000 158.4440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.2440 0.0000 158.4440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 158.2440 0.0000 158.4440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 158.2440 0.0000 158.4440 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[114]

  PIN I[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.9270 0.0000 159.1270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.9270 0.0000 159.1270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.9270 0.0000 159.1270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 158.9270 0.0000 159.1270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 158.9270 0.0000 159.1270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[115]

  PIN O[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 160.9800 0.0000 161.1800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.9800 0.0000 161.1800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.9800 0.0000 161.1800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 160.9800 0.0000 161.1800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 160.9800 0.0000 161.1800 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[116]

  PIN O[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 159.6120 0.0000 159.8120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 159.6120 0.0000 159.8120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 159.6120 0.0000 159.8120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 159.6120 0.0000 159.8120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 159.6120 0.0000 159.8120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[115]

  PIN I[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 160.2950 0.0000 160.4950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.2950 0.0000 160.4950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.2950 0.0000 160.4950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 160.2950 0.0000 160.4950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 160.2950 0.0000 160.4950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[116]

  PIN I[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 161.6630 0.0000 161.8630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.6630 0.0000 161.8630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.6630 0.0000 161.8630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 161.6630 0.0000 161.8630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 161.6630 0.0000 161.8630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[117]

  PIN O[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 162.3480 0.0000 162.5480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 162.3480 0.0000 162.5480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 162.3480 0.0000 162.5480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 162.3480 0.0000 162.5480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 162.3480 0.0000 162.5480 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[117]

  PIN I[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 163.0310 0.0000 163.2310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 163.0310 0.0000 163.2310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 163.0310 0.0000 163.2310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 163.0310 0.0000 163.2310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 163.0310 0.0000 163.2310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[118]

  PIN O[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 163.7160 0.0000 163.9160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 163.7160 0.0000 163.9160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 163.7160 0.0000 163.9160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 163.7160 0.0000 163.9160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 163.7160 0.0000 163.9160 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[118]

  PIN I[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 164.3990 0.0000 164.5990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.3990 0.0000 164.5990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.3990 0.0000 164.5990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 164.3990 0.0000 164.5990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 164.3990 0.0000 164.5990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[119]

  PIN O[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 165.0840 0.0000 165.2840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.0840 0.0000 165.2840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.0840 0.0000 165.2840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 165.0840 0.0000 165.2840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 165.0840 0.0000 165.2840 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 25.3008 LAYER M4 ;
    ANTENNADIFFAREA 1843.297 LAYER M5 ;
    ANTENNADIFFAREA 1843.297 LAYER M6 ;
    ANTENNADIFFAREA 1843.297 LAYER M7 ;
    ANTENNADIFFAREA 1843.297 LAYER M8 ;
    ANTENNADIFFAREA 1843.297 LAYER M9 ;
    ANTENNADIFFAREA 1843.297 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 2.6394 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 402.6647 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 402.6647 LAYER M4 ;
    ANTENNAMAXAREACAR 165.8826 LAYER M4 ;
    ANTENNAGATEAREA 11.0823 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 18045.2 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 18045.2 LAYER M5 ;
    ANTENNAMAXAREACAR 1794.895 LAYER M5 ;
    ANTENNAGATEAREA 11.0823 LAYER M6 ;
    ANTENNAGATEAREA 11.0823 LAYER M7 ;
    ANTENNAGATEAREA 11.0823 LAYER M8 ;
    ANTENNAGATEAREA 11.0823 LAYER M9 ;
    ANTENNAGATEAREA 11.0823 LAYER MRDL ;
  END O[119]

  PIN I[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 165.7670 0.0000 165.9670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.7670 0.0000 165.9670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.7670 0.0000 165.9670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 165.7670 0.0000 165.9670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 165.7670 0.0000 165.9670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[120]

  PIN O[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 166.4520 0.0000 166.6520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 166.4520 0.0000 166.6520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 166.4520 0.0000 166.6520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 166.4520 0.0000 166.6520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 166.4520 0.0000 166.6520 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[120]

  PIN I[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 167.1350 0.0000 167.3350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.1350 0.0000 167.3350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.1350 0.0000 167.3350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 167.1350 0.0000 167.3350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 167.1350 0.0000 167.3350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[121]

  PIN O[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 167.8200 0.0000 168.0200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.8200 0.0000 168.0200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.8200 0.0000 168.0200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 167.8200 0.0000 168.0200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 167.8200 0.0000 168.0200 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[121]

  PIN I[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 168.5030 0.0000 168.7030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.5030 0.0000 168.7030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.5030 0.0000 168.7030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 168.5030 0.0000 168.7030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 168.5030 0.0000 168.7030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[122]

  PIN O[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 169.1880 0.0000 169.3880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.1880 0.0000 169.3880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.1880 0.0000 169.3880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 169.1880 0.0000 169.3880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 169.1880 0.0000 169.3880 0.2000 ;
    END
    ANTENNADIFFAREA 1.091992 LAYER M3 ;
    ANTENNADIFFAREA 1.091992 LAYER M4 ;
    ANTENNADIFFAREA 1.091992 LAYER M5 ;
    ANTENNADIFFAREA 1.091992 LAYER M6 ;
    ANTENNADIFFAREA 1.091992 LAYER M7 ;
    ANTENNADIFFAREA 1.091992 LAYER M8 ;
    ANTENNADIFFAREA 1.091992 LAYER M9 ;
    ANTENNADIFFAREA 1.091992 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 2.079404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.079404 LAYER M3 ;
    ANTENNAMAXAREACAR 100.2675 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END O[122]

  PIN I[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 143.8790 0.0000 144.0790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.8790 0.0000 144.0790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.8790 0.0000 144.0790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 143.8790 0.0000 144.0790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 143.8790 0.0000 144.0790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[104]

  PIN O[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 144.5640 0.0000 144.7640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.5640 0.0000 144.7640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.5640 0.0000 144.7640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 144.5640 0.0000 144.7640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 144.5640 0.0000 144.7640 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[104]

  PIN I[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 145.2470 0.0000 145.4470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.2470 0.0000 145.4470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.2470 0.0000 145.4470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 145.2470 0.0000 145.4470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 145.2470 0.0000 145.4470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[105]

  PIN O[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 145.9320 0.0000 146.1320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.9320 0.0000 146.1320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.9320 0.0000 146.1320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 145.9320 0.0000 146.1320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 145.9320 0.0000 146.1320 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[105]

  PIN I[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 146.6150 0.0000 146.8150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.6150 0.0000 146.8150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.6150 0.0000 146.8150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 146.6150 0.0000 146.8150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 146.6150 0.0000 146.8150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[106]

  PIN O[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 147.3000 0.0000 147.5000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.3000 0.0000 147.5000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.3000 0.0000 147.5000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 147.3000 0.0000 147.5000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 147.3000 0.0000 147.5000 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[106]

  PIN I[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 147.9830 0.0000 148.1830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.9830 0.0000 148.1830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.9830 0.0000 148.1830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 147.9830 0.0000 148.1830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 147.9830 0.0000 148.1830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[107]

  PIN O[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 148.6680 0.0000 148.8680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.6680 0.0000 148.8680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.6680 0.0000 148.8680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 148.6680 0.0000 148.8680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 148.6680 0.0000 148.8680 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[107]

  PIN I[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 149.3510 0.0000 149.5510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.3510 0.0000 149.5510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.3510 0.0000 149.5510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 149.3510 0.0000 149.5510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 149.3510 0.0000 149.5510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[108]

  PIN O[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.0360 0.0000 150.2360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.0360 0.0000 150.2360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.0360 0.0000 150.2360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.0360 0.0000 150.2360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.0360 0.0000 150.2360 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[108]

  PIN I[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 150.7190 0.0000 150.9190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.7190 0.0000 150.9190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.7190 0.0000 150.9190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 150.7190 0.0000 150.9190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 150.7190 0.0000 150.9190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[109]

  PIN O[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 151.4040 0.0000 151.6040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 151.4040 0.0000 151.6040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 151.4040 0.0000 151.6040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 151.4040 0.0000 151.6040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 151.4040 0.0000 151.6040 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[109]

  PIN I[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 152.0870 0.0000 152.2870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.0870 0.0000 152.2870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.0870 0.0000 152.2870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 152.0870 0.0000 152.2870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 152.0870 0.0000 152.2870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[110]

  PIN O[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 152.7720 0.0000 152.9720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.7720 0.0000 152.9720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.7720 0.0000 152.9720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 152.7720 0.0000 152.9720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 152.7720 0.0000 152.9720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[110]

  PIN I[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 153.4550 0.0000 153.6550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.4550 0.0000 153.6550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.4550 0.0000 153.6550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 153.4550 0.0000 153.6550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 153.4550 0.0000 153.6550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[111]

  PIN O[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.1400 0.0000 154.3400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.1400 0.0000 154.3400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.1400 0.0000 154.3400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.1400 0.0000 154.3400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.1400 0.0000 154.3400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[111]

  PIN I[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 154.8230 0.0000 155.0230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.8230 0.0000 155.0230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.8230 0.0000 155.0230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 154.8230 0.0000 155.0230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 154.8230 0.0000 155.0230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[112]

  PIN O[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 155.5080 0.0000 155.7080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 155.5080 0.0000 155.7080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 155.5080 0.0000 155.7080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 155.5080 0.0000 155.7080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 155.5080 0.0000 155.7080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[112]

  PIN I[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 156.1910 0.0000 156.3910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.1910 0.0000 156.3910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.1910 0.0000 156.3910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 156.1910 0.0000 156.3910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 156.1910 0.0000 156.3910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[113]

  PIN I[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 131.5670 0.0000 131.7670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.5670 0.0000 131.7670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.5670 0.0000 131.7670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 131.5670 0.0000 131.7670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 131.5670 0.0000 131.7670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[95]

  PIN O[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.2520 0.0000 132.4520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.2520 0.0000 132.4520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.2520 0.0000 132.4520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.2520 0.0000 132.4520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.2520 0.0000 132.4520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[95]

  PIN I[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 132.9350 0.0000 133.1350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.9350 0.0000 133.1350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.9350 0.0000 133.1350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 132.9350 0.0000 133.1350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 132.9350 0.0000 133.1350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[96]

  PIN O[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 133.6200 0.0000 133.8200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.6200 0.0000 133.8200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.6200 0.0000 133.8200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 133.6200 0.0000 133.8200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 133.6200 0.0000 133.8200 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[96]

  PIN I[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 134.3030 0.0000 134.5030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.3030 0.0000 134.5030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.3030 0.0000 134.5030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.3030 0.0000 134.5030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 134.3030 0.0000 134.5030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[97]

  PIN O[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 134.9880 0.0000 135.1880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.9880 0.0000 135.1880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.9880 0.0000 135.1880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 134.9880 0.0000 135.1880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 134.9880 0.0000 135.1880 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[97]

  PIN I[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 130.1990 0.0000 130.3990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.1990 0.0000 130.3990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.1990 0.0000 130.3990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 130.1990 0.0000 130.3990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 130.1990 0.0000 130.3990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[94]

  PIN I[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 135.6710 0.0000 135.8710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 135.6710 0.0000 135.8710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 135.6710 0.0000 135.8710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 135.6710 0.0000 135.8710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 135.6710 0.0000 135.8710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[98]

  PIN I[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 137.0390 0.0000 137.2390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.0390 0.0000 137.2390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.0390 0.0000 137.2390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 137.0390 0.0000 137.2390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 137.0390 0.0000 137.2390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[99]

  PIN O[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 137.7240 0.0000 137.9240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.7240 0.0000 137.9240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.7240 0.0000 137.9240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 137.7240 0.0000 137.9240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 137.7240 0.0000 137.9240 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[99]

  PIN I[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 138.4070 0.0000 138.6070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.4070 0.0000 138.6070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.4070 0.0000 138.6070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 138.4070 0.0000 138.6070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 138.4070 0.0000 138.6070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[100]

  PIN O[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 139.0920 0.0000 139.2920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.0920 0.0000 139.2920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.0920 0.0000 139.2920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 139.0920 0.0000 139.2920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 139.0920 0.0000 139.2920 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[100]

  PIN I[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 139.7750 0.0000 139.9750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.7750 0.0000 139.9750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.7750 0.0000 139.9750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 139.7750 0.0000 139.9750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 139.7750 0.0000 139.9750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[101]

  PIN O[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 140.4600 0.0000 140.6600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 140.4600 0.0000 140.6600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 140.4600 0.0000 140.6600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 140.4600 0.0000 140.6600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 140.4600 0.0000 140.6600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[101]

  PIN I[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 141.1430 0.0000 141.3430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.1430 0.0000 141.3430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.1430 0.0000 141.3430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 141.1430 0.0000 141.3430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 141.1430 0.0000 141.3430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[102]

  PIN O[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 141.8280 0.0000 142.0280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.8280 0.0000 142.0280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.8280 0.0000 142.0280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 141.8280 0.0000 142.0280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 141.8280 0.0000 142.0280 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[102]

  PIN I[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 142.5110 0.0000 142.7110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.5110 0.0000 142.7110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.5110 0.0000 142.7110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 142.5110 0.0000 142.7110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 142.5110 0.0000 142.7110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[103]

  PIN O[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 143.1960 0.0000 143.3960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.1960 0.0000 143.3960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.1960 0.0000 143.3960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 143.1960 0.0000 143.3960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 143.1960 0.0000 143.3960 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[103]

  PIN O[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 118.5720 0.0000 118.7720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.5720 0.0000 118.7720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.5720 0.0000 118.7720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 118.5720 0.0000 118.7720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 118.5720 0.0000 118.7720 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[85]

  PIN I[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 119.2550 0.0000 119.4550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.2550 0.0000 119.4550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.2550 0.0000 119.4550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.2550 0.0000 119.4550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.2550 0.0000 119.4550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[86]

  PIN O[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 119.9400 0.0000 120.1400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.9400 0.0000 120.1400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.9400 0.0000 120.1400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 119.9400 0.0000 120.1400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 119.9400 0.0000 120.1400 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[86]

  PIN I[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 120.6230 0.0000 120.8230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.6230 0.0000 120.8230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.6230 0.0000 120.8230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 120.6230 0.0000 120.8230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 120.6230 0.0000 120.8230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[87]

  PIN O[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 121.3080 0.0000 121.5080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.3080 0.0000 121.5080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.3080 0.0000 121.5080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 121.3080 0.0000 121.5080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.3080 0.0000 121.5080 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.274264 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[87]

  PIN I[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 121.9910 0.0000 122.1910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.9910 0.0000 122.1910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.9910 0.0000 122.1910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 121.9910 0.0000 122.1910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 121.9910 0.0000 122.1910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28374 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28374 LAYER M3 ;
    ANTENNAMAXAREACAR 62.37874 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.59367 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 76.80813 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[88]
  OBS
    LAYER M1 ;
      RECT 196.7220 115.6650 197.5220 115.8550 ;
      RECT 0.0000 0.0000 1.0070 0.8000 ;
      RECT 196.0210 131.1910 197.5220 133.0430 ;
      RECT 0.0000 0.8000 197.5220 9.2200 ;
      RECT 177.5010 0.0000 197.5220 9.2200 ;
      RECT 177.5010 0.0000 197.5220 0.8000 ;
      RECT 0.0000 117.2550 197.5220 123.0850 ;
      RECT 0.0000 114.2650 196.7220 117.2550 ;
      RECT 0.0000 108.4230 197.5220 114.2650 ;
      RECT 0.0000 105.4450 196.7220 108.4230 ;
      RECT 0.0000 99.5070 197.5220 105.4450 ;
      RECT 0.0000 98.1070 196.7220 99.5070 ;
      RECT 0.0000 18.0900 197.5220 98.1070 ;
      RECT 0.0000 16.2280 196.7220 18.0900 ;
      RECT 0.0000 10.6200 197.5220 16.2280 ;
      RECT 0.0000 9.2200 196.7210 10.6200 ;
      RECT 0.0000 134.4430 197.5220 140.7440 ;
      RECT 0.0000 124.4850 196.7280 140.7440 ;
      RECT 0.0000 10.6200 196.7220 140.7440 ;
      RECT 0.0000 10.6200 196.7220 140.7440 ;
      RECT 0.0000 10.6200 196.7220 140.7440 ;
      RECT 0.0000 10.6200 196.7220 140.7440 ;
      RECT 0.0000 10.6200 196.7220 140.7440 ;
      RECT 0.0000 0.8000 196.7210 140.7440 ;
      RECT 0.0000 129.4480 196.7280 134.4430 ;
      RECT 0.0000 124.4850 197.5220 129.4480 ;
      RECT 0.0000 123.0850 196.7220 124.4850 ;
      RECT 196.7220 106.8450 197.5220 107.0230 ;
    LAYER PO ;
      RECT 0.0000 0.0000 197.5220 140.7440 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 197.5220 140.7440 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 197.5220 140.7440 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 197.5220 140.7440 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 197.5220 140.7440 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 197.5220 140.7440 ;
    LAYER M5 ;
      RECT 0.0000 139.7440 0.2120 140.7440 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 0.0000 0.0000 0.9070 0.9010 ;
      RECT 197.2110 139.7440 197.5220 140.7440 ;
      RECT 0.0000 0.9000 2.2750 0.9010 ;
      RECT 0.0000 0.9000 2.2750 2.4010 ;
      RECT 196.0210 131.2910 197.5220 132.9430 ;
      RECT 177.6010 0.0000 197.5220 0.9000 ;
      RECT 0.0000 0.9010 197.5220 9.1200 ;
      RECT 3.8750 0.9000 65.2030 0.9010 ;
      RECT 66.8030 0.9000 128.1310 0.9010 ;
      RECT 129.7310 0.9000 197.5220 9.1200 ;
      RECT 129.7310 0.9000 197.5220 0.9010 ;
      RECT 0.0000 117.3550 197.5220 122.9850 ;
      RECT 0.0000 114.1650 196.6220 117.3550 ;
      RECT 0.0000 108.5230 197.5220 114.1650 ;
      RECT 0.0000 105.3450 196.6220 108.5230 ;
      RECT 0.0000 99.6070 197.5220 105.3450 ;
      RECT 0.0000 98.0070 196.6220 99.6070 ;
      RECT 0.0000 18.1900 197.5220 98.0070 ;
      RECT 0.0000 16.1280 196.6220 18.1900 ;
      RECT 0.0000 10.7200 197.5220 16.1280 ;
      RECT 0.0000 9.1200 196.6210 10.7200 ;
      RECT 0.0000 134.5430 197.5220 139.7440 ;
      RECT 0.0000 124.5850 196.6280 139.7440 ;
      RECT 0.0000 10.7200 196.6220 139.7440 ;
      RECT 0.0000 10.7200 196.6220 139.7440 ;
      RECT 0.0000 10.7200 196.6220 139.7440 ;
      RECT 0.0000 10.7200 196.6220 139.7440 ;
      RECT 0.0000 10.7200 196.6220 139.7440 ;
      RECT 0.0000 0.9010 196.6210 139.7440 ;
      RECT 0.0000 129.3480 196.6280 134.5430 ;
      RECT 0.0000 124.5850 197.5220 129.3480 ;
      RECT 0.0000 122.9850 196.6220 124.5850 ;
      RECT 3.8750 0.9000 65.2030 139.7440 ;
      RECT 66.8030 0.9000 128.1310 139.7440 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 0.0000 0.0000 0.9070 0.9010 ;
      RECT 0.0000 0.9000 2.2750 2.4010 ;
      RECT 196.0210 131.2910 197.5220 132.9430 ;
      RECT 177.6010 0.0000 197.5220 0.9000 ;
      RECT 0.0000 0.9010 197.5220 9.1200 ;
      RECT 3.8750 0.9000 65.2030 0.9010 ;
      RECT 66.8030 0.9000 128.1310 0.9010 ;
      RECT 129.7310 0.9000 197.5220 9.1200 ;
      RECT 129.7310 0.9000 197.5220 0.9010 ;
      RECT 0.0000 117.3550 197.5220 122.9850 ;
      RECT 0.0000 114.1650 196.6220 117.3550 ;
      RECT 0.0000 108.5230 197.5220 114.1650 ;
      RECT 0.0000 105.3450 196.6220 108.5230 ;
      RECT 0.0000 99.6070 197.5220 105.3450 ;
      RECT 0.0000 98.0070 196.6220 99.6070 ;
      RECT 0.0000 18.1900 197.5220 98.0070 ;
      RECT 0.0000 16.1280 196.6220 18.1900 ;
      RECT 0.0000 10.7200 197.5220 16.1280 ;
      RECT 0.0000 9.1200 196.6210 10.7200 ;
      RECT 0.0000 134.5430 197.5220 140.7440 ;
      RECT 0.0000 124.5850 196.6280 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 0.9010 196.6210 140.7440 ;
      RECT 0.0000 129.3480 196.6280 134.5430 ;
      RECT 0.0000 124.5850 197.5220 129.3480 ;
      RECT 0.0000 122.9850 196.6220 124.5850 ;
      RECT 3.8750 0.9000 65.2030 140.7440 ;
      RECT 66.8030 0.9000 128.1310 140.7440 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 196.0210 131.2910 197.5220 132.9430 ;
      RECT 0.0000 0.9000 197.5220 9.1200 ;
      RECT 177.6010 0.0000 197.5220 9.1200 ;
      RECT 177.6010 0.0000 197.5220 0.9000 ;
      RECT 0.0000 117.3550 197.5220 122.9850 ;
      RECT 0.0000 114.1650 196.6220 117.3550 ;
      RECT 0.0000 108.5230 197.5220 114.1650 ;
      RECT 0.0000 105.3450 196.6220 108.5230 ;
      RECT 0.0000 99.6070 197.5220 105.3450 ;
      RECT 0.0000 98.0070 196.6220 99.6070 ;
      RECT 0.0000 18.1900 197.5220 98.0070 ;
      RECT 0.0000 16.1280 196.6220 18.1900 ;
      RECT 0.0000 10.7200 197.5220 16.1280 ;
      RECT 0.0000 9.1200 196.6210 10.7200 ;
      RECT 0.0000 134.5430 197.5220 140.7440 ;
      RECT 0.0000 124.5850 196.6280 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 0.9000 196.6210 140.7440 ;
      RECT 0.0000 129.3480 196.6280 134.5430 ;
      RECT 0.0000 124.5850 197.5220 129.3480 ;
      RECT 0.0000 122.9850 196.6220 124.5850 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 196.0210 131.2910 197.5220 132.9430 ;
      RECT 0.0000 0.9000 197.5220 9.1200 ;
      RECT 177.6010 0.0000 197.5220 9.1200 ;
      RECT 177.6010 0.0000 197.5220 0.9000 ;
      RECT 0.0000 117.3550 197.5220 122.9850 ;
      RECT 0.0000 114.1650 196.6220 117.3550 ;
      RECT 0.0000 108.5230 197.5220 114.1650 ;
      RECT 0.0000 105.3450 196.6220 108.5230 ;
      RECT 0.0000 99.6070 197.5220 105.3450 ;
      RECT 0.0000 98.0070 196.6220 99.6070 ;
      RECT 0.0000 18.1900 197.5220 98.0070 ;
      RECT 0.0000 16.1280 196.6220 18.1900 ;
      RECT 0.0000 10.7200 197.5220 16.1280 ;
      RECT 0.0000 9.1200 196.6210 10.7200 ;
      RECT 0.0000 134.5430 197.5220 140.7440 ;
      RECT 0.0000 124.5850 196.6280 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 10.7200 196.6220 140.7440 ;
      RECT 0.0000 0.9000 196.6210 140.7440 ;
      RECT 0.0000 129.3480 196.6280 134.5430 ;
      RECT 0.0000 124.5850 197.5220 129.3480 ;
      RECT 0.0000 122.9850 196.6220 124.5850 ;
  END
END SRAMLP1RW64x128

MACRO SRAMLP1RW128x8
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 33.302 BY 240.241 ;
  SYMMETRY X Y R90 ;

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2600 0.0000 2.4600 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[0]

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3420 0.0000 4.5420 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[1]

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0780 0.0000 7.2780 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[4]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0070 0.0000 5.2070 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[1]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6370 0.0000 3.8370 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[7]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9740 0.0000 3.1740 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[7]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 185.3330 33.3020 185.5330 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 185.3330 33.3020 185.5330 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 185.3330 33.3020 185.5330 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 185.3330 33.3020 185.5330 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 185.3330 33.3020 185.5330 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END A[4]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 16.8990 33.3020 17.0990 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 16.8990 33.3020 17.0990 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 16.8990 33.3020 17.0990 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 16.8990 33.3020 17.0990 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 16.8990 33.3020 17.0990 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15058 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15058 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15058 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.15058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15058 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.423229 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.423229 LAYER M4 ;
    ANTENNAMAXAREACAR 14.25845 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 18.36679 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1080 205.8110 33.3020 206.0110 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1080 205.8110 33.3020 206.0110 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1080 205.8110 33.3020 206.0110 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1080 205.8110 33.3020 206.0110 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1080 205.8110 33.3020 206.0110 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END SD

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6060 0.0000 1.8060 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[0]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 178.1120 33.3020 178.3120 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 178.1120 33.3020 178.3120 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 178.1120 33.3020 178.3120 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 178.1120 33.3020 178.3120 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 178.1120 33.3020 178.3120 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END A[5]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1080 209.3130 33.3020 209.5130 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1080 209.3130 33.3020 209.5130 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1080 209.3130 33.3020 209.5130 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1080 209.3130 33.3020 209.5130 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1080 209.3130 33.3020 209.5130 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.280905 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.280905 LAYER M1 ;
    ANTENNAGATEAREA 0.0366 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END LS

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 186.9310 33.3020 187.1310 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 186.9310 33.3020 187.1310 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 186.9310 33.3020 187.1310 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 186.9310 33.3020 187.1310 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 186.9310 33.3020 187.1310 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 30.8757 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 440.2544 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 440.2544 LAYER M1 ;
    ANTENNAGATEAREA 40.4202 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 695.2174 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 695.2174 LAYER M2 ;
    ANTENNAMAXAREACAR 29.36906 LAYER M2 ;
    ANTENNAGATEAREA 40.4202 LAYER M3 ;
    ANTENNAGATEAREA 40.4202 LAYER M4 ;
    ANTENNAGATEAREA 40.4202 LAYER M5 ;
    ANTENNAGATEAREA 40.4202 LAYER M6 ;
    ANTENNAGATEAREA 40.4202 LAYER M7 ;
    ANTENNAGATEAREA 40.4202 LAYER M8 ;
    ANTENNAGATEAREA 40.4202 LAYER M9 ;
    ANTENNAGATEAREA 40.4202 LAYER MRDL ;
  END A[3]

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1080 206.1910 33.3020 206.3910 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1080 206.1910 33.3020 206.3910 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1080 206.1910 33.3020 206.3910 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1080 206.1910 33.3020 206.3910 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1080 206.1910 33.3020 206.3910 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END DS

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 194.1530 33.3020 194.3530 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 194.1530 33.3020 194.3530 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 194.1530 33.3020 194.3530 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 194.1530 33.3020 194.3530 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 194.1530 33.3020 194.3530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END A[2]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 176.5150 33.3020 176.7150 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 176.5150 33.3020 176.7150 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 176.5150 33.3020 176.7150 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 176.5150 33.3020 176.7150 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 176.5150 33.3020 176.7150 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
    ANTENNAGATEAREA 48.3468 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 115.243 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.243 LAYER M3 ;
    ANTENNAMAXAREACAR 10.01618 LAYER M3 ;
    ANTENNAGATEAREA 48.3468 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 729.7753 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 729.7753 LAYER M4 ;
    ANTENNAMAXAREACAR 48.93695 LAYER M4 ;
    ANTENNAGATEAREA 52.6326 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 5154.164 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 5154.164 LAYER M5 ;
    ANTENNAMAXAREACAR 215.51 LAYER M5 ;
    ANTENNAGATEAREA 52.6326 LAYER M6 ;
    ANTENNAGATEAREA 52.6326 LAYER M7 ;
    ANTENNAGATEAREA 52.6326 LAYER M8 ;
    ANTENNAGATEAREA 52.6326 LAYER M9 ;
    ANTENNAGATEAREA 52.6326 LAYER MRDL ;
  END A[6]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 195.7530 33.3020 195.9530 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 195.7530 33.3020 195.9530 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 195.7530 33.3020 195.9530 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 195.7530 33.3020 195.9530 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 195.7530 33.3020 195.9530 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END A[1]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 9.8900 33.3020 10.0900 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 9.8900 33.3020 10.0900 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 9.8900 33.3020 10.0900 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 9.8900 33.3020 10.0900 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 9.8900 33.3020 10.0900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.56544 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.56544 LAYER M2 ;
    ANTENNAMAXAREACAR 11.75319 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 12.79006 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 13.82686 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 14.86359 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 202.9700 33.3020 203.1700 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 202.9700 33.3020 203.1700 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 202.9700 33.3020 203.1700 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 202.9700 33.3020 203.1700 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 202.9700 33.3020 203.1700 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1507 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1507 LAYER M2 ;
  END A[0]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.1020 17.3590 33.3020 17.5590 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.1020 17.3590 33.3020 17.5590 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.1020 17.3590 33.3020 17.5590 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.1020 17.3590 33.3020 17.5590 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.1020 17.3590 33.3020 17.5590 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.15058 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15058 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.15058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15058 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.15058 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15058 LAYER M3 ;
    ANTENNAGATEAREA 0.0342 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.30412 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.30412 LAYER M4 ;
    ANTENNAMAXAREACAR 13.40876 LAYER M4 ;
    ANTENNAGATEAREA 0.0342 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1504 LAYER M5 ;
    ANTENNAMAXAREACAR 17.80553 LAYER M5 ;
    ANTENNAGATEAREA 0.0342 LAYER M6 ;
    ANTENNAGATEAREA 0.0342 LAYER M7 ;
    ANTENNAGATEAREA 0.0342 LAYER M8 ;
    ANTENNAGATEAREA 0.0342 LAYER M9 ;
    ANTENNAGATEAREA 0.0342 LAYER MRDL ;
  END CE

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 3.7020 239.9410 4.0020 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.6010 239.9410 4.9010 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.4010 239.9410 24.7000 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.3010 239.9410 25.6000 240.2410 ;
    END
  END VDDL

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8140 0.0000 10.0140 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[3]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5500 0.0000 12.7500 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1434 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.91606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.91606 LAYER M2 ;
    ANTENNAMAXAREACAR 7.35416 LAYER M2 ;
    ANTENNAGATEAREA 0.1434 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAMAXAREACAR 8.410858 LAYER M3 ;
    ANTENNAGATEAREA 0.1434 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 9.467485 LAYER M4 ;
    ANTENNAGATEAREA 0.1434 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 10.52404 LAYER M5 ;
    ANTENNAGATEAREA 0.1434 LAYER M6 ;
    ANTENNAGATEAREA 0.1434 LAYER M7 ;
    ANTENNAGATEAREA 0.1434 LAYER M8 ;
    ANTENNAGATEAREA 0.1434 LAYER M9 ;
    ANTENNAGATEAREA 0.1434 LAYER MRDL ;
  END OEB

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1820 0.0000 11.3820 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[5]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1120 0.0000 9.3120 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[2]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 29.8010 239.9410 30.1000 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.7010 239.9410 31.0010 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.0010 239.9410 1.3020 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.1020 239.9410 0.4010 240.2410 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 4.1510 239.9410 4.4520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.0510 239.9410 14.3510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.4510 239.9410 10.7510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.3520 239.9410 2.6510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.8520 239.9410 16.1520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.7510 239.9410 17.0500 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.9510 239.9410 15.2510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.6520 239.9410 17.9530 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.8520 239.9410 7.1520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.3520 239.9410 11.6520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.1520 239.9410 13.4530 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.2510 239.9410 12.5500 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.7510 239.9410 8.0500 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.5510 239.9410 9.8510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.6520 239.9410 8.9530 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.1510 239.9410 31.4510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.5520 239.9410 27.8520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.9520 239.9410 24.2520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.3520 239.9410 20.6520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.5510 239.9410 18.8510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.0520 239.9410 32.3520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.2510 239.9410 30.5510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.3510 239.9410 29.6510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.4510 239.9410 28.7510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.6510 239.9410 26.9510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.7510 239.9410 26.0510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.8510 239.9410 25.1510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.0510 239.9410 23.3510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.1510 239.9410 22.4510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.2510 239.9410 21.5510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.4510 239.9410 19.7510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.4520 239.9410 1.7510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.5520 239.9410 0.8520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.0510 239.9410 5.3510 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.2510 239.9410 3.5520 240.2410 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.9510 239.9410 6.2510 240.2410 ;
    END
  END VSS

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8520 0.0000 12.0520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[5]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.4820 0.0000 10.6820 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[3]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4460 0.0000 8.6460 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[2]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7300 0.0000 7.9300 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277608 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[4]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7100 0.0000 5.9100 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.021 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.28812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.28812 LAYER M3 ;
    ANTENNAMAXAREACAR 62.58731 LAYER M3 ;
    ANTENNAGATEAREA 0.021 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 69.80223 LAYER M4 ;
    ANTENNAGATEAREA 0.021 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 77.01667 LAYER M5 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ;
    ANTENNAGATEAREA 0.021 LAYER M7 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ;
    ANTENNAGATEAREA 0.021 LAYER MRDL ;
  END I[6]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3760 0.0000 6.5760 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.277728 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[6]
  OBS
    LAYER M1 ;
      RECT 13.3500 0.0000 33.3020 9.2900 ;
      RECT 13.3500 0.0000 33.3020 0.8000 ;
      RECT 0.0000 210.1130 33.3020 240.2410 ;
      RECT 0.0000 203.7700 32.5080 240.2410 ;
      RECT 0.0000 0.8000 32.5020 240.2410 ;
      RECT 0.0000 0.8000 32.5020 240.2410 ;
      RECT 0.0000 0.8000 32.5020 240.2410 ;
      RECT 0.0000 0.8000 32.5020 240.2410 ;
      RECT 0.0000 0.8000 32.5020 240.2410 ;
      RECT 0.0000 0.8000 32.5020 240.2410 ;
      RECT 0.0000 203.7700 32.5080 210.1130 ;
      RECT 0.0000 202.3700 32.5020 203.7700 ;
      RECT 32.5020 194.9530 33.3020 195.1530 ;
      RECT 32.5020 177.3150 33.3020 177.5120 ;
      RECT 32.5020 186.1330 33.3020 186.3310 ;
      RECT 0.0000 0.0000 1.0060 0.8000 ;
      RECT 32.5080 203.7700 33.3020 205.2110 ;
      RECT 31.8010 206.9910 33.3020 208.7130 ;
      RECT 0.0000 196.5530 33.3020 202.3700 ;
      RECT 0.0000 193.5530 32.5020 196.5530 ;
      RECT 0.0000 187.7310 33.3020 193.5530 ;
      RECT 0.0000 184.7330 32.5020 187.7310 ;
      RECT 0.0000 178.9120 33.3020 184.7330 ;
      RECT 0.0000 175.9150 32.5020 178.9120 ;
      RECT 0.0000 18.1590 33.3020 175.9150 ;
      RECT 0.0000 16.2990 32.5020 18.1590 ;
      RECT 0.0000 10.6900 33.3020 16.2990 ;
      RECT 0.0000 9.2900 32.5020 10.6900 ;
      RECT 0.0000 0.8000 33.3020 9.2900 ;
    LAYER PO ;
      RECT 0.0000 0.0000 33.3020 240.2410 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 33.3020 240.2410 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 33.3020 240.2410 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 33.3020 240.2410 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 33.3020 240.2410 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 33.3020 240.2410 ;
    LAYER M5 ;
      RECT 33.0520 239.2410 33.3020 240.2410 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.8010 207.0910 33.3020 208.6130 ;
      RECT 32.4080 203.8700 33.3020 205.1110 ;
      RECT 0.0000 196.6530 33.3020 202.2700 ;
      RECT 0.0000 193.4530 32.4020 196.6530 ;
      RECT 0.0000 187.8310 33.3020 193.4530 ;
      RECT 0.0000 184.6330 32.4020 187.8310 ;
      RECT 0.0000 179.0120 33.3020 184.6330 ;
      RECT 0.0000 175.8150 32.4020 179.0120 ;
      RECT 0.0000 18.2590 33.3020 175.8150 ;
      RECT 0.0000 16.1990 32.4020 18.2590 ;
      RECT 0.0000 10.7900 33.3020 16.1990 ;
      RECT 0.0000 9.1900 32.4020 10.7900 ;
      RECT 0.0000 0.9000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 0.9000 ;
      RECT 0.0000 210.2130 33.3020 239.2410 ;
      RECT 0.0000 203.8700 32.4080 239.2410 ;
      RECT 0.0000 0.9000 32.4020 239.2410 ;
      RECT 0.0000 0.9000 32.4020 239.2410 ;
      RECT 0.0000 0.9000 32.4020 239.2410 ;
      RECT 0.0000 0.9000 32.4020 239.2410 ;
      RECT 0.0000 0.9000 32.4020 239.2410 ;
      RECT 0.0000 0.9000 32.4020 239.2410 ;
      RECT 0.0000 203.8700 32.4080 210.2130 ;
      RECT 0.0000 202.2700 32.4020 203.8700 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.8010 207.0910 33.3020 208.6130 ;
      RECT 32.4080 203.8700 33.3020 205.1110 ;
      RECT 0.0000 196.6530 33.3020 202.2700 ;
      RECT 0.0000 193.4530 32.4020 196.6530 ;
      RECT 0.0000 187.8310 33.3020 193.4530 ;
      RECT 0.0000 184.6330 32.4020 187.8310 ;
      RECT 0.0000 179.0120 33.3020 184.6330 ;
      RECT 0.0000 175.8150 32.4020 179.0120 ;
      RECT 0.0000 18.2590 33.3020 175.8150 ;
      RECT 0.0000 16.1990 32.4020 18.2590 ;
      RECT 0.0000 10.7900 33.3020 16.1990 ;
      RECT 0.0000 9.1900 32.4020 10.7900 ;
      RECT 0.0000 0.9000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 0.9000 ;
      RECT 0.0000 210.2130 33.3020 240.2410 ;
      RECT 0.0000 203.8700 32.4080 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 203.8700 32.4080 210.2130 ;
      RECT 0.0000 202.2700 32.4020 203.8700 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 31.8010 207.0910 33.3020 208.6130 ;
      RECT 32.4080 203.8700 33.3020 205.1110 ;
      RECT 0.0000 196.6530 33.3020 202.2700 ;
      RECT 0.0000 193.4530 32.4020 196.6530 ;
      RECT 0.0000 187.8310 33.3020 193.4530 ;
      RECT 0.0000 184.6330 32.4020 187.8310 ;
      RECT 0.0000 179.0120 33.3020 184.6330 ;
      RECT 0.0000 175.8150 32.4020 179.0120 ;
      RECT 0.0000 18.2590 33.3020 175.8150 ;
      RECT 0.0000 16.1990 32.4020 18.2590 ;
      RECT 0.0000 10.7900 33.3020 16.1990 ;
      RECT 0.0000 9.1900 32.4020 10.7900 ;
      RECT 0.0000 0.9000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 0.9000 ;
      RECT 0.0000 210.2130 33.3020 240.2410 ;
      RECT 0.0000 203.8700 32.4080 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 203.8700 32.4080 210.2130 ;
      RECT 0.0000 202.2700 32.4020 203.8700 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 0.9060 0.9000 ;
      RECT 32.4080 203.8700 33.3020 205.1110 ;
      RECT 31.8010 207.0910 33.3020 208.6130 ;
      RECT 0.0000 196.6530 33.3020 202.2700 ;
      RECT 0.0000 193.4530 32.4020 196.6530 ;
      RECT 0.0000 187.8310 33.3020 193.4530 ;
      RECT 0.0000 184.6330 32.4020 187.8310 ;
      RECT 0.0000 179.0120 33.3020 184.6330 ;
      RECT 0.0000 175.8150 32.4020 179.0120 ;
      RECT 0.0000 18.2590 33.3020 175.8150 ;
      RECT 0.0000 16.1990 32.4020 18.2590 ;
      RECT 0.0000 10.7900 33.3020 16.1990 ;
      RECT 0.0000 9.1900 32.4020 10.7900 ;
      RECT 0.0000 0.9000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 9.1900 ;
      RECT 13.4500 0.0000 33.3020 0.9000 ;
      RECT 0.0000 210.2130 33.3020 240.2410 ;
      RECT 0.0000 203.8700 32.4080 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 0.9000 32.4020 240.2410 ;
      RECT 0.0000 203.8700 32.4080 210.2130 ;
      RECT 0.0000 202.2700 32.4020 203.8700 ;
  END
END SRAMLP1RW128x8

MACRO SRAMLP1RW128x46
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 93.899 BY 240.379 ;
  SYMMETRY X Y R90 ;

  PIN I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 60.4310 0.0000 60.6310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[10]

  PIN O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.7480 0.0000 59.9480 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[11]

  PIN O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 21.4440 0.0000 21.6440 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[14]

  PIN I[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.1270 0.0000 22.3270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[40]

  PIN I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.9670 0.0000 29.1670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[9]

  PIN O[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 28.2840 0.0000 28.4840 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[32]

  PIN I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 34.4390 0.0000 34.6390 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[7]

  PIN O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 47.4360 0.0000 47.6360 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[20]

  PIN I[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 42.6470 0.0000 42.8470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[44]

  PIN O[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.9640 0.0000 42.1640 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[43]

  PIN O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.7560 0.0000 33.9560 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[8]

  PIN I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.1190 0.0000 48.3190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[28]

  PIN I[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 27.5990 0.0000 27.7990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[32]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 0.7910 240.0790 1.0910 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.6900 240.0790 1.9890 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.1850 240.0790 87.4840 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.0850 240.0790 88.3840 240.3790 ;
    END
  END VDD

  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 186.8560 93.8990 187.0560 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 186.8560 93.8990 187.0560 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 186.8560 93.8990 187.0560 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 186.8560 93.8990 187.0560 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 186.8560 93.8990 187.0560 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.5068 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5068 LAYER M3 ;
    ANTENNAMAXAREACAR 33.48762 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.62749 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 41.76708 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[3]

  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 185.5660 93.8990 185.7660 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 185.5660 93.8990 185.7660 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 185.5660 93.8990 185.7660 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 185.5660 93.8990 185.7660 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 185.5660 93.8990 185.7660 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.52924 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52924 LAYER M3 ;
    ANTENNAMAXAREACAR 34.09665 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 38.23648 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.37604 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[4]

  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 178.0400 93.8990 178.2400 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 178.0400 93.8990 178.2400 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 178.0400 93.8990 178.2400 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 178.0400 93.8990 178.2400 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 178.0400 93.8990 178.2400 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.5263 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5263 LAYER M3 ;
    ANTENNAMAXAREACAR 33.75951 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.89935 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.03893 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[5]

  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 176.4500 93.8990 176.6500 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 176.4500 93.8990 176.6500 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 176.4500 93.8990 176.6500 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 176.4500 93.8990 176.6500 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 176.4500 93.8990 176.6500 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.5263 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5263 LAYER M3 ;
    ANTENNAMAXAREACAR 33.75814 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.89799 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.03757 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[6]

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 17.2900 93.8990 17.4900 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 17.2900 93.8990 17.4900 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 17.2900 93.8990 17.4900 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 17.2900 93.8990 17.4900 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 17.2900 93.8990 17.4900 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0576 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 3.00598 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.00598 LAYER M4 ;
    ANTENNAMAXAREACAR 65.57839 LAYER M4 ;
    ANTENNAGATEAREA 0.0576 LAYER M5 ;
    ANTENNAGATEAREA 0.0576 LAYER M6 ;
    ANTENNAGATEAREA 0.0576 LAYER M7 ;
    ANTENNAGATEAREA 0.0576 LAYER M8 ;
    ANTENNAGATEAREA 0.0576 LAYER M9 ;
    ANTENNAGATEAREA 0.0576 LAYER MRDL ;
  END CE

  PIN I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.6070 0.0000 1.8070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 24.6465 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 535.551 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 535.551 LAYER M3 ;
    ANTENNAMAXAREACAR 2340.119 LAYER M3 ;
    ANTENNAGATEAREA 24.6465 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 2839.849 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2839.849 LAYER M4 ;
    ANTENNAMAXAREACAR 2455.343 LAYER M4 ;
    ANTENNAGATEAREA 77.3409 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 14308.96 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 14308.96 LAYER M5 ;
    ANTENNAMAXAREACAR 264.1412 LAYER M5 ;
    ANTENNAGATEAREA 77.3409 LAYER M6 ;
    ANTENNAGATEAREA 77.3409 LAYER M7 ;
    ANTENNAGATEAREA 77.3409 LAYER M8 ;
    ANTENNAGATEAREA 77.3409 LAYER M9 ;
    ANTENNAGATEAREA 77.3409 LAYER MRDL ;
  END I[4]

  PIN CSB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 16.8280 93.8990 17.0280 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 16.8280 93.8990 17.0280 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 16.8280 93.8990 17.0280 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 16.8280 93.8990 17.0280 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 16.8280 93.8990 17.0280 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.947029 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.947029 LAYER M4 ;
    ANTENNAMAXAREACAR 29.13688 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 33.27704 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END CSB

  PIN I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.7990 0.0000 61.9990 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[15]

  PIN O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 6.3960 0.0000 6.5960 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[18]

  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 229.6290 93.8990 229.8290 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 229.6290 93.8990 229.8290 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 229.6290 93.8990 229.8290 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 229.6290 93.8990 229.8290 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 229.6290 93.8990 229.8290 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.2256 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.146276 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.146276 LAYER M2 ;
    ANTENNAMAXAREACAR 9.885359 LAYER M2 ;
    ANTENNAGATEAREA 36.5436 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 18.53301 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.53301 LAYER M3 ;
    ANTENNAMAXAREACAR 16.19187 LAYER M3 ;
    ANTENNAGATEAREA 36.5436 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 308.068 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 308.068 LAYER M4 ;
    ANTENNAMAXAREACAR 26.43102 LAYER M4 ;
    ANTENNAGATEAREA 36.5436 LAYER M5 ;
    ANTENNAGATEAREA 36.5436 LAYER M6 ;
    ANTENNAGATEAREA 36.5436 LAYER M7 ;
    ANTENNAGATEAREA 36.5436 LAYER M8 ;
    ANTENNAGATEAREA 36.5436 LAYER M9 ;
    ANTENNAGATEAREA 36.5436 LAYER MRDL ;
  END SD

  PIN VDDL
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 2.5910 240.0790 2.8920 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.4900 240.0790 3.7900 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.3860 240.0790 85.6860 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.2850 240.0790 86.5840 240.3790 ;
    END
  END VDDL

  PIN DS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 230.3920 93.8990 230.5920 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 230.3920 93.8990 230.5920 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 230.3920 93.8990 230.5920 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 230.3920 93.8990 230.5920 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 230.3920 93.8990 230.5920 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
  END DS

  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 202.9060 93.8990 203.1060 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 202.9060 93.8990 203.1060 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 202.9060 93.8990 203.1060 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 202.9060 93.8990 203.1060 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 202.9060 93.8990 203.1060 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.5263 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5263 LAYER M3 ;
    ANTENNAMAXAREACAR 33.73901 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.87886 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.01844 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[0]

  PIN LS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 233.5490 93.8990 233.7490 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 233.5490 93.8990 233.7490 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 233.5490 93.8990 233.7490 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 233.5490 93.8990 233.7490 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 233.5490 93.8990 233.7490 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAGATEAREA 0.0366 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.593101 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.593101 LAYER M1 ;
    ANTENNAGATEAREA 23.3598 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 30.1058 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1058 LAYER M2 ;
    ANTENNAMAXAREACAR 5.792699 LAYER M2 ;
    ANTENNAGATEAREA 23.3598 LAYER M3 ;
    ANTENNAGATEAREA 23.3598 LAYER M4 ;
    ANTENNAGATEAREA 23.3598 LAYER M5 ;
    ANTENNAGATEAREA 23.3598 LAYER M6 ;
    ANTENNAGATEAREA 23.3598 LAYER M7 ;
    ANTENNAGATEAREA 23.3598 LAYER M8 ;
    ANTENNAGATEAREA 23.3598 LAYER M9 ;
    ANTENNAGATEAREA 23.3598 LAYER MRDL ;
  END LS

  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 194.0860 93.8990 194.2860 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 194.0860 93.8990 194.2860 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 194.0860 93.8990 194.2860 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 194.0860 93.8990 194.2860 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 194.0860 93.8990 194.2860 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.5263 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5263 LAYER M3 ;
    ANTENNAMAXAREACAR 33.72125 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 37.86111 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.00069 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[2]

  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 195.6760 93.8990 195.8760 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 195.6760 93.8990 195.8760 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 195.6760 93.8990 195.8760 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 195.6760 93.8990 195.8760 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 195.6760 93.8990 195.8760 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAGATEAREA 0.0366 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.7519 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7519 LAYER M3 ;
    ANTENNAMAXAREACAR 34.70462 LAYER M3 ;
    ANTENNAGATEAREA 0.0366 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 38.84441 LAYER M4 ;
    ANTENNAGATEAREA 0.0366 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 42.98392 LAYER M5 ;
    ANTENNAGATEAREA 0.0366 LAYER M6 ;
    ANTENNAGATEAREA 0.0366 LAYER M7 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ;
    ANTENNAGATEAREA 0.0366 LAYER M9 ;
    ANTENNAGATEAREA 0.0366 LAYER MRDL ;
  END A[1]

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 90.3340 240.0780 90.6340 240.3780 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.2360 240.0780 91.5360 240.3780 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.4350 240.0780 89.7350 240.3780 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.1350 240.0780 92.4350 240.3780 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.3410 240.0790 0.6420 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 1.2400 240.0790 1.5400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.9400 240.0790 4.2390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.5340 240.0790 88.8340 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.4400 240.0790 8.7400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 2.1400 240.0790 2.4400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.7400 240.0790 6.0400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.2400 240.0790 10.5400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.3400 240.0790 9.6400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.8400 240.0790 14.1400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.9400 240.0790 13.2400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.7410 240.0790 15.0410 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.6350 240.0790 87.9350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.5410 240.0790 7.8410 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.1410 240.0790 11.4410 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.2390 240.0790 19.5390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.0400 240.0790 12.3400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.5400 240.0790 16.8400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.6400 240.0790 15.9400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.4390 240.0790 17.7390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.1390 240.0790 20.4390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.0390 240.0790 21.3380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.3400 240.0790 18.6400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.7380 240.0790 24.0390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.6380 240.0790 24.9380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.8380 240.0790 23.1390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.4390 240.0790 26.7390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.1380 240.0790 29.4380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.9390 240.0790 22.2380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.5380 240.0790 25.8380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.3380 240.0790 27.6370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.2390 240.0790 28.5400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.0380 240.0790 30.3380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.9390 240.0790 31.2390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.7390 240.0790 33.0400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.8380 240.0790 32.1370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.5380 240.0790 34.8380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.6380 240.0790 33.9380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.1380 240.0790 38.4380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.4390 240.0790 35.7390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.0380 240.0790 39.3380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.2390 240.0790 37.5400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.6380 240.0790 42.9380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.3380 240.0790 36.6370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.8380 240.0790 41.1380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.5390 240.0790 43.8390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.7380 240.0790 42.0380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.9380 240.0790 49.2380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.0380 240.0790 48.3380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.9390 240.0790 40.2390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.3380 240.0790 45.6380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.4380 240.0790 44.7380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.2380 240.0790 46.5380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.5360 240.0790 52.8360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.4360 240.0790 53.7350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.1390 240.0790 47.4390 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.8370 240.0790 50.1370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.7380 240.0790 51.0380 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.6370 240.0790 51.9370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.1350 240.0790 56.4360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.9350 240.0790 58.2350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.2350 240.0790 55.5360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.3360 240.0790 54.6350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.4350 240.0790 62.7350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.0350 240.0790 57.3350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.8360 240.0790 59.1360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.5350 240.0790 61.8350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.3360 240.0790 63.6360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.7350 240.0790 60.0340 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.9350 240.0790 67.2350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.6360 240.0790 60.9370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.0350 240.0790 66.3350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.2350 240.0790 64.5340 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.8360 240.0790 68.1360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.4350 240.0790 71.7350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.3360 240.0790 72.6360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.1360 240.0790 65.4370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.7350 240.0790 69.0340 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.6360 240.0790 69.9370 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.5350 240.0790 70.8350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.8350 240.0790 77.1350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.0350 240.0790 75.3350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.7350 240.0790 78.0350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.2350 240.0790 73.5350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.9360 240.0790 76.2360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.1350 240.0790 74.4350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.3350 240.0790 81.6350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.4350 240.0790 80.7350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.2340 240.0790 82.5340 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.5360 240.0790 79.8360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.7350 240.0790 87.0350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.6350 240.0790 78.9350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.0340 240.0790 84.3340 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.0410 240.0790 3.3410 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.8360 240.0790 86.1360 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.6400 240.0790 6.9400 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.1350 240.0790 83.4350 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.8410 240.0790 5.1420 240.3790 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.9350 240.0790 85.2350 240.3790 ;
    END
    ANTENNAPARTIALMETALAREA 71.8344 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 71.8344 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 71.8344 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 71.8344 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 71.8338 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 71.8338 LAYER M5 ;
  END VSS

  PIN I[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.9590 0.0000 55.1590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[38]

  PIN I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.7510 0.0000 46.9510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[20]

  PIN O[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.1800 0.0000 24.3800 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[37]

  PIN I[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 56.3270 0.0000 56.5270 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[33]

  PIN O[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.0120 0.0000 57.2120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[33]

  PIN I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.1830 0.0000 11.3830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[22]

  PIN O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 58.3800 0.0000 58.5800 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[12]

  PIN I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 59.0630 0.0000 59.2630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[11]

  PIN O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 10.5000 0.0000 10.7000 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[21]

  PIN I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 4.3430 0.0000 4.5430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[16]

  PIN I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 57.6950 0.0000 57.8950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[12]

  PIN I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.1670 0.0000 63.3670 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[30]

  PIN O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 63.8520 0.0000 64.0520 0.2000 ;
    END
    ANTENNADIFFAREA 0.11118 LAYER M3 ;
    ANTENNADIFFAREA 0.11118 LAYER M4 ;
    ANTENNADIFFAREA 0.11118 LAYER M5 ;
    ANTENNADIFFAREA 0.11118 LAYER M6 ;
    ANTENNADIFFAREA 0.11118 LAYER M7 ;
    ANTENNADIFFAREA 0.11118 LAYER M8 ;
    ANTENNADIFFAREA 0.11118 LAYER M9 ;
    ANTENNADIFFAREA 0.11118 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.280384 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.280384 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
  END O[30]

  PIN O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 62.4840 0.0000 62.6840 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[15]

  PIN OEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 64.5250 0.0000 64.7250 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.5250 0.0000 64.7250 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.5250 0.0000 64.7250 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 64.5250 0.0000 64.7250 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 64.5250 0.0000 64.7250 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 1.0956 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 8.21008 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.21008 LAYER M2 ;
    ANTENNAMAXAREACAR 38.91342 LAYER M2 ;
    ANTENNAGATEAREA 1.0956 LAYER M3 ;
    ANTENNAGATEAREA 1.0956 LAYER M4 ;
    ANTENNAGATEAREA 1.0956 LAYER M5 ;
    ANTENNAGATEAREA 1.0956 LAYER M6 ;
    ANTENNAGATEAREA 1.0956 LAYER M7 ;
    ANTENNAGATEAREA 1.0956 LAYER M8 ;
    ANTENNAGATEAREA 1.0956 LAYER M9 ;
    ANTENNAGATEAREA 1.0956 LAYER MRDL ;
  END OEB

  PIN O[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 55.6440 0.0000 55.8440 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[38]

  PIN O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.6520 0.0000 29.8520 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[9]

  PIN O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 14.6040 0.0000 14.8040 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[24]

  PIN O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.7000 0.0000 44.9000 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[0]

  PIN I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.2870 0.0000 15.4870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[25]

  PIN O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 40.5960 0.0000 40.7960 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[3]

  PIN I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 44.0150 0.0000 44.2150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[0]

  PIN O[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 25.5480 0.0000 25.7480 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[34]

  PIN I[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 24.8630 0.0000 25.0630 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[34]

  PIN O[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 46.0680 0.0000 46.2680 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[45]

  PIN I[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 45.3830 0.0000 45.5830 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[45]

  PIN I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 12.5510 0.0000 12.7510 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[23]

  PIN O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 11.8680 0.0000 12.0680 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[22]

  PIN O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.1320 0.0000 9.3320 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[29]

  PIN I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.9190 0.0000 14.1190 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[24]

  PIN O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 13.2360 0.0000 13.4360 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[23]

  PIN I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.8150 0.0000 10.0150 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[21]

  PIN O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 51.5400 0.0000 51.7400 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[19]

  PIN I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.2230 0.0000 52.4230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[17]

  PIN O[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 54.2760 0.0000 54.4760 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[42]

  PIN O[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 43.3320 0.0000 43.5320 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[44]

  PIN O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.0280 0.0000 5.2280 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[16]

  PIN O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 3.6600 0.0000 3.8600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[2]

  PIN I[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 41.2790 0.0000 41.4790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[43]

  PIN I[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.7030 0.0000 31.9030 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[36]

  PIN I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.7590 0.0000 20.9590 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[14]

  PIN O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 20.0760 0.0000 20.2760 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[13]

  PIN O[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 31.0200 0.0000 31.2200 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[35]

  PIN O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.7080 0.0000 18.9080 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[27]

  PIN O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 15.9720 0.0000 16.1720 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[25]

  PIN I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 19.3910 0.0000 19.5910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[13]

  PIN I[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 16.6550 0.0000 16.8550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[41]

  PIN I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.1750 0.0000 37.3750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[6]

  PIN I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.2310 0.0000 26.4310 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[31]

  PIN O[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 36.4920 0.0000 36.6920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[39]

  PIN I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 33.0710 0.0000 33.2710 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[8]

  PIN O[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 32.3880 0.0000 32.5880 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[36]

  PIN I[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 30.3350 0.0000 30.5350 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[35]

  PIN O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 26.9160 0.0000 27.1160 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[31]

  PIN I[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.8070 0.0000 36.0070 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[39]

  PIN O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 35.1240 0.0000 35.3240 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[7]

  PIN I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 49.4870 0.0000 49.6870 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[26]

  PIN O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.1720 0.0000 50.3720 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[26]

  PIN I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 50.8550 0.0000 51.0550 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[19]

  PIN O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 48.8040 0.0000 49.0040 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[28]

  PIN I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 38.5430 0.0000 38.7430 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[5]

  PIN O[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 22.8120 0.0000 23.0120 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[40]

  PIN I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 18.0230 0.0000 18.2230 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[27]

  PIN O[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 17.3400 0.0000 17.5400 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[41]

  PIN O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 37.8600 0.0000 38.0600 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[6]

  PIN I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.9110 0.0000 40.1110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[3]

  PIN I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.9750 0.0010 3.1750 0.2010 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.9750 0.0010 3.1750 0.2010 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.9750 0.0000 3.1750 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[2]

  PIN I[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 23.4950 0.0000 23.6950 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[37]

  PIN O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 39.2280 0.0000 39.4280 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[5]

  PIN O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 2.2920 0.0000 2.4920 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[4]

  PIN I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 8.4470 0.0000 8.6470 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[29]

  PIN O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.7640 0.0000 7.9640 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[1]

  PIN WEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 93.6990 9.8200 93.8990 10.0200 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.6990 9.8200 93.8990 10.0200 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.6990 9.8200 93.8990 10.0200 ;
    END
    PORT
      LAYER M2 ;
        RECT 93.6990 9.8200 93.8990 10.0200 ;
    END
    PORT
      LAYER M1 ;
        RECT 93.6990 9.8200 93.8990 10.0200 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAGATEAREA 0.1461 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 2.08222 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.08222 LAYER M2 ;
    ANTENNAMAXAREACAR 15.29036 LAYER M2 ;
    ANTENNAGATEAREA 0.1461 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.1525 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1525 LAYER M3 ;
    ANTENNAMAXAREACAR 16.33316 LAYER M3 ;
    ANTENNAGATEAREA 0.1461 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M4 ;
    ANTENNAMAXAREACAR 17.36973 LAYER M4 ;
    ANTENNAGATEAREA 0.1461 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M5 ;
    ANTENNAMAXAREACAR 18.40623 LAYER M5 ;
    ANTENNAGATEAREA 0.1461 LAYER M6 ;
    ANTENNAGATEAREA 0.1461 LAYER M7 ;
    ANTENNAGATEAREA 0.1461 LAYER M8 ;
    ANTENNAGATEAREA 0.1461 LAYER M9 ;
    ANTENNAGATEAREA 0.1461 LAYER MRDL ;
  END WEB

  PIN I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 7.0790 0.0000 7.2790 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[1]

  PIN I[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 53.5910 0.0000 53.7910 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[42]

  PIN O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 52.9080 0.0000 53.1080 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[17]

  PIN I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.7110 0.0000 5.9110 0.2000 ;
    END
    ANTENNADIFFAREA 0.6 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END I[18]

  PIN O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M2 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    PORT
      LAYER M1 ;
        RECT 61.1160 0.0000 61.3160 0.2000 ;
    END
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0.1516 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1516 LAYER M2 ;
  END O[10]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
      RECT 0.0000 229.0290 93.0990 234.3490 ;
      RECT 0.0000 203.7060 93.8990 229.0290 ;
      RECT 0.0000 202.3060 93.0990 203.7060 ;
      RECT 0.0000 196.4760 93.8990 202.3060 ;
      RECT 0.0000 193.4860 93.0990 196.4760 ;
      RECT 0.0000 187.6560 93.8990 193.4860 ;
      RECT 0.0000 184.9660 93.0990 187.6560 ;
      RECT 0.0000 178.8400 93.8990 184.9660 ;
      RECT 0.0000 175.8500 93.0990 178.8400 ;
      RECT 0.0000 18.0900 93.8990 175.8500 ;
      RECT 0.0000 16.2280 93.0990 18.0900 ;
      RECT 0.0000 10.6200 93.8990 16.2280 ;
      RECT 0.0000 9.2200 93.0990 10.6200 ;
      RECT 0.0000 0.8000 93.8990 9.2200 ;
      RECT 65.3250 0.0000 93.8990 9.2200 ;
      RECT 65.3250 0.0000 93.8990 0.8000 ;
      RECT 93.0990 177.2500 93.8990 177.4400 ;
      RECT 93.0990 194.8860 93.8990 195.0760 ;
      RECT 0.0000 0.0000 1.0070 0.8000 ;
      RECT 92.3980 231.1920 93.8990 232.9490 ;
      RECT 0.0000 234.3490 93.8990 240.3790 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
      RECT 0.0000 0.8000 93.0990 240.3790 ;
    LAYER PO ;
      RECT 0.0000 0.0000 93.8990 240.3790 ;
    LAYER MRDL ;
      RECT 0.0000 0.0000 93.8990 240.3790 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 93.8990 240.3790 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 93.8990 240.3790 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 93.8990 240.3790 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 93.8990 240.3790 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 0.9070 0.9010 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 93.1350 239.3780 93.8990 240.3790 ;
      RECT 0.0000 0.9000 2.2750 0.9010 ;
      RECT 0.0000 0.9000 2.2750 2.4010 ;
      RECT 92.3980 231.2920 93.8990 232.8490 ;
      RECT 65.4250 0.0000 93.8990 0.9000 ;
      RECT 0.0000 239.3780 88.7350 239.3790 ;
      RECT 0.0000 0.9010 88.7350 239.3790 ;
      RECT 0.0000 234.4490 93.8990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 0.9010 92.9990 239.3780 ;
      RECT 0.0000 228.9290 92.9990 234.4490 ;
      RECT 0.0000 203.8060 93.8990 228.9290 ;
      RECT 0.0000 202.2060 92.9990 203.8060 ;
      RECT 0.0000 196.5760 93.8990 202.2060 ;
      RECT 0.0000 193.3860 92.9990 196.5760 ;
      RECT 0.0000 187.7560 93.8990 193.3860 ;
      RECT 0.0000 184.8660 92.9990 187.7560 ;
      RECT 0.0000 178.9400 93.8990 184.8660 ;
      RECT 0.0000 175.7500 92.9990 178.9400 ;
      RECT 0.0000 18.1900 93.8990 175.7500 ;
      RECT 0.0000 16.1280 92.9990 18.1900 ;
      RECT 0.0000 10.7200 93.8990 16.1280 ;
      RECT 0.0000 9.1200 92.9990 10.7200 ;
      RECT 0.0000 0.9010 93.8990 9.1200 ;
      RECT 3.8750 0.9000 93.8990 9.1200 ;
      RECT 3.8750 0.9000 93.8990 0.9010 ;
      RECT 65.4250 0.0000 93.8990 9.1200 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 0.0000 0.9000 2.2750 2.4010 ;
      RECT 92.3980 231.2920 93.8990 232.8490 ;
      RECT 65.4250 0.0000 93.8990 0.9000 ;
      RECT 0.0000 234.4490 93.8990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 0.9010 92.9990 240.3790 ;
      RECT 0.0000 228.9290 92.9990 234.4490 ;
      RECT 0.0000 203.8060 93.8990 228.9290 ;
      RECT 0.0000 202.2060 92.9990 203.8060 ;
      RECT 0.0000 196.5760 93.8990 202.2060 ;
      RECT 0.0000 193.3860 92.9990 196.5760 ;
      RECT 0.0000 187.7560 93.8990 193.3860 ;
      RECT 0.0000 184.8660 92.9990 187.7560 ;
      RECT 0.0000 178.9400 93.8990 184.8660 ;
      RECT 0.0000 175.7500 92.9990 178.9400 ;
      RECT 0.0000 18.1900 93.8990 175.7500 ;
      RECT 0.0000 16.1280 92.9990 18.1900 ;
      RECT 0.0000 10.7200 93.8990 16.1280 ;
      RECT 0.0000 9.1200 92.9990 10.7200 ;
      RECT 0.0000 0.9010 93.8990 9.1200 ;
      RECT 3.8750 0.9000 93.8990 9.1200 ;
      RECT 3.8750 0.9000 93.8990 0.9010 ;
      RECT 65.4250 0.0000 93.8990 9.1200 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 92.3980 231.2920 93.8990 232.8490 ;
      RECT 0.0000 234.4490 93.8990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 228.9290 92.9990 234.4490 ;
      RECT 0.0000 203.8060 93.8990 228.9290 ;
      RECT 0.0000 202.2060 92.9990 203.8060 ;
      RECT 0.0000 196.5760 93.8990 202.2060 ;
      RECT 0.0000 193.3860 92.9990 196.5760 ;
      RECT 0.0000 187.7560 93.8990 193.3860 ;
      RECT 0.0000 184.8660 92.9990 187.7560 ;
      RECT 0.0000 178.9400 93.8990 184.8660 ;
      RECT 0.0000 175.7500 92.9990 178.9400 ;
      RECT 0.0000 18.1900 93.8990 175.7500 ;
      RECT 0.0000 16.1280 92.9990 18.1900 ;
      RECT 0.0000 10.7200 93.8990 16.1280 ;
      RECT 0.0000 9.1200 92.9990 10.7200 ;
      RECT 0.0000 0.9000 93.8990 9.1200 ;
      RECT 65.4250 0.0000 93.8990 9.1200 ;
      RECT 65.4250 0.0000 93.8990 0.9000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 0.9070 0.9000 ;
      RECT 92.3980 231.2920 93.8990 232.8490 ;
      RECT 0.0000 234.4490 93.8990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 0.9000 92.9990 240.3790 ;
      RECT 0.0000 228.9290 92.9990 234.4490 ;
      RECT 0.0000 203.8060 93.8990 228.9290 ;
      RECT 0.0000 202.2060 92.9990 203.8060 ;
      RECT 0.0000 196.5760 93.8990 202.2060 ;
      RECT 0.0000 193.3860 92.9990 196.5760 ;
      RECT 0.0000 187.7560 93.8990 193.3860 ;
      RECT 0.0000 184.8660 92.9990 187.7560 ;
      RECT 0.0000 178.9400 93.8990 184.8660 ;
      RECT 0.0000 175.7500 92.9990 178.9400 ;
      RECT 0.0000 18.1900 93.8990 175.7500 ;
      RECT 0.0000 16.1280 92.9990 18.1900 ;
      RECT 0.0000 10.7200 93.8990 16.1280 ;
      RECT 0.0000 9.1200 92.9990 10.7200 ;
      RECT 0.0000 0.9000 93.8990 9.1200 ;
      RECT 65.4250 0.0000 93.8990 9.1200 ;
      RECT 65.4250 0.0000 93.8990 0.9000 ;
  END
END SRAMLP1RW128x46
  
END LIBRARY
